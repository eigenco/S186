// vi: ft=systemverilog
//`ifndef MICROCODE_ROM_PATH
//`define MICROCODE_ROM_PATH "."
//`endif

//`default_nettype none
module Microcode(input logic clk,
                 input logic reset,
                 input logic nmi_pulse,
                 input logic intr,
                 output logic inta,
                 output logic irq_to_mdr,
                 output logic start_interrupt,
                 output logic do_escape_fault,
                 output logic starting_instruction,
                 input logic stall,
                 input logic divide_error,
                 input logic rm_is_reg,
                 input logic [2:0] modrm_reg,
                 input logic int_enabled,
                 input logic zf,
                 input logic tf,
                 output logic [15:0] microcode_immediate,
                 output logic [8:0] update_flags,
                 output logic modrm_start,
                 output logic use_microcode_immediate,
                 output logic [7:0] opcode,
                 input logic jump_taken,
                 input logic rb_zero,
                 output logic lock,
                 output logic multibit_shift,
                 output logic is_hlt,
                 output logic next_microinstruction,
                 // Microinstruction fields.
                 output logic [1:0] a_sel,
                 output logic [5:0] alu_op,
                 output logic [2:0] b_sel,
                 output logic ext_int_yield,
                 output logic io,
                 output logic load_ip,
                 output logic mar_wr_sel,
                 output logic mar_write,
                 output logic mdr_write,
                 output logic mem_read,
                 output logic mem_write,
                 output logic next_instruction,
                 output logic ra_modrm_rm_reg,
                 output logic [2:0] ra_sel,
                 output logic rb_cl,
                 output logic [2:0] rd_sel,
                 output logic [1:0] rd_sel_source,
                 output logic [1:0] reg_wr_source,
                 output logic [1:0] segment,
                 output logic segment_force,
                 output logic segment_wr_en,
                 output logic tmp_wr_en,
                 output logic tmp_wr_sel,
                 output logic width,
                 output logic reg_wr_en,
                 // Fifo Read Port.
                 output logic fifo_rd_en,
                 // verilator lint_off UNUSED
                 input Instruction next_instruction_value,
                 output Instruction cur_instruction,
                 // verilator lint_on UNUSED
                 input logic fifo_empty,
                 input logic fifo_resetting,
                 output logic loop_next,
                 input logic loop_done,
                 // Debug
                 output logic debug_stopped,
                 input logic debug_seize,
                 input logic [7:0] debug_addr,
                 input logic debug_run);

localparam num_instructions = 1196;
localparam addr_bits = 11;
localparam reset_address = 11'h129;
localparam nmi_address = 11'h12a;
localparam irq_address = 11'h12b;
localparam single_step_address = 11'h12c;
localparam divide_error_address = 11'h101;
localparam next_instruction_address = 11'h100;
localparam modrm_wait_address = 11'h12e;
localparam bad_opcode_address = 11'h12f;
localparam debug_wait_address = 11'h102;
localparam do_int_address = 11'h12d;

typedef struct packed {
    logic [10:0] next;
    logic [1:0] a_sel;
    logic [5:0] alu_op;
    logic [2:0] b_sel;
    logic ext_int_inhibit;
    logic ext_int_yield;
    logic [3:0] immediate;
    logic io;
    logic [3:0] jump_type;
    logic load_ip;
    logic mar_wr_sel;
    logic mar_write;
    logic mdr_write;
    logic mem_read;
    logic mem_write;
    logic next_instruction;
    logic ra_modrm_rm_reg;
    logic [2:0] ra_sel;
    logic rb_cl;
    logic [2:0] rd_sel;
    logic [1:0] rd_sel_source;
    logic [1:0] reg_wr_source;
    logic [1:0] segment;
    logic segment_force;
    logic segment_wr_en;
    logic tmp_wr_en;
    logic tmp_wr_sel;
    logic [3:0] update_flags;
    logic [1:0] width;
} microcode_instruction;

microcode_instruction mem[num_instructions];
microcode_instruction current;
reg [addr_bits-1:0] addr;
reg [addr_bits-1:0] next_addr;
reg [addr_bits-1:0] jump_target;
assign use_microcode_immediate = |current.immediate;
assign opcode = cur_instruction.opcode;

initial
begin
mem[0] = 64'b0010100010100000000000000000000010010000100000000000110000000010;
mem[1] = 64'b0010100010100000000000000000000010010000100000000000110000000010;
mem[2] = 64'b0010100100000000000000000000000010010000100000000000110000000010;
mem[3] = 64'b0010100100000000000000000000000010010000100000000000110000000010;
mem[4] = 64'b0010100101100000000000000000000000000000000000000000000000000010;
mem[5] = 64'b0010100101100000000000000000000000000000000000000000000000000010;
mem[6] = 64'b0110010111000000000000000000000000000000000000000000001000000000;
mem[7] = 64'b0101111111100000000000000000000000000000010000000000000000000000;
mem[8] = 64'b0101110100000000000000000000000010010000100000000000110000000010;
mem[9] = 64'b0101110100000000000000000000000010010000100000000000110000000010;
mem[10] = 64'b0101110101100000000000000000000010010000100000000000110000000010;
mem[11] = 64'b0101110101100000000000000000000010010000100000000000110000000010;
mem[12] = 64'b0101110111000000000000000000000000000000000000000000000000000010;
mem[13] = 64'b0101110111000000000000000000000000000000000000000000000000000010;
mem[14] = 64'b0110010111000000000000000000000000000000000000000000011000000000;
mem[15] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[16] = 64'b0010011011000000000000000000000010010000100000000000110000000010;
mem[17] = 64'b0010011011000000000000000000000010010000100000000000110000000010;
mem[18] = 64'b0010011100100000000000000000000010010000100000000000110000000010;
mem[19] = 64'b0010011100100000000000000000000010010000100000000000110000000010;
mem[20] = 64'b0010011110000000000000000000000000000000000000000000000000000010;
mem[21] = 64'b0010011110000000000000000000000000000000000000000000000000000010;
mem[22] = 64'b0110010111000000000000000000000000000000000000000000101000000000;
mem[23] = 64'b0110000001000000000000000000000000000000010000000000000000000000;
mem[24] = 64'b0111010101000000000000000000000010010000100000000000110000000010;
mem[25] = 64'b0111010101000000000000000000000010010000100000000000110000000010;
mem[26] = 64'b0111010110100000000000000000000010010000100000000000110000000010;
mem[27] = 64'b0111010110100000000000000000000010010000100000000000110000000010;
mem[28] = 64'b0111011000000000000000000000000000000000000000000000000000000010;
mem[29] = 64'b0111011000000000000000000000000000000000000000000000000000000010;
mem[30] = 64'b0110010111000000000000000000000000000000000000000000111000000000;
mem[31] = 64'b0110000010100000000000000000000000000000010000000000000000000000;
mem[32] = 64'b0010101010000000000000000000000010010000100000000000110000000010;
mem[33] = 64'b0010101010000000000000000000000010010000100000000000110000000010;
mem[34] = 64'b0010101011100000000000000000000010010000100000000000110000000010;
mem[35] = 64'b0010101011100000000000000000000010010000100000000000110000000010;
mem[36] = 64'b0010101101000000000000000000000000000000000000000000000000000010;
mem[37] = 64'b0010101101000000000000000000000000000000000000000000000000000010;
mem[38] = 64'b0000010011100000000000000000000000000001000000000000000000000000;
mem[39] = 64'b0010110110100000000000000000000000000000000000000000000000000000;
mem[40] = 64'b0111111001000000000000000000000010010000100000000000110000000010;
mem[41] = 64'b0111111001000000000000000000000010010000100000000000110000000010;
mem[42] = 64'b0111111010100000000000000000000010010000100000000000110000000010;
mem[43] = 64'b0111111010100000000000000000000010010000100000000000110000000010;
mem[44] = 64'b0111111100000000000000000000000000000000000000000000000000000010;
mem[45] = 64'b0111111100000000000000000000000000000000000000000000000000000010;
mem[46] = 64'b0000010111100000000000000000000000000001000000000000000000000000;
mem[47] = 64'b0010110111000000000000000000000000000000000000000000000000000000;
mem[48] = 64'b1000010101100000000000000000000010010000100000000000110000000010;
mem[49] = 64'b1000010101100000000000000000000010010000100000000000110000000010;
mem[50] = 64'b1000010111000000000000000000000010010000100000000000110000000010;
mem[51] = 64'b1000010111000000000000000000000010010000100000000000110000000010;
mem[52] = 64'b1000011000100000000000000000000000000000000000000000000000000010;
mem[53] = 64'b1000011000100000000000000000000000000000000000000000000000000010;
mem[54] = 64'b0000011011100000000000000000000000000001000000000000000000000000;
mem[55] = 64'b0010011000000000000000000000000000000000000000000000000000000000;
mem[56] = 64'b0011000110000000000000000000000010010000100000000000110000000010;
mem[57] = 64'b0011000110000000000000000000000010010000100000000000110000000010;
mem[58] = 64'b0011000111100000000000000000000010010000100000000000110000000010;
mem[59] = 64'b0011000111100000000000000000000010010000100000000000110000000010;
mem[60] = 64'b0011001001000000000000000000000000000000000000000000000000000010;
mem[61] = 64'b0011001001000000000000000000000000000000000000000000000000000010;
mem[62] = 64'b0000011111100000000000000000000000000001000000000000000000000000;
mem[63] = 64'b0010011010100000000000000000000000000000000000000000000000000000;
mem[64] = 64'b0011111011000000000000000000000000000000000000000000000000000000;
mem[65] = 64'b0011111011100000000000000000000000000000000100000000000000000000;
mem[66] = 64'b0011111100000000000000000000000000000000001000000000000000000000;
mem[67] = 64'b0011111100100000000000000000000000000000001100000000000000000000;
mem[68] = 64'b0011111101000000000000000000000000000000010000000000000000000000;
mem[69] = 64'b0011111101100000000000000000000000000000010100000000000000000000;
mem[70] = 64'b0011111110000000000000000000000000000000011000000000000000000000;
mem[71] = 64'b0011111110100000000000000000000000000000011100000000000000000000;
mem[72] = 64'b0011111111000000000000000000000000000000000000000000000000000000;
mem[73] = 64'b0011111111100000000000000000000000000000000100000000000000000000;
mem[74] = 64'b0100000000000000000000000000000000000000001000000000000000000000;
mem[75] = 64'b0100000000100000000000000000000000000000001100000000000000000000;
mem[76] = 64'b0100000001000000000000000000000000000000010000000000000000000000;
mem[77] = 64'b0100000001100000000000000000000000000000010100000000000000000000;
mem[78] = 64'b0100000010000000000000000000000000000000011000000000000000000000;
mem[79] = 64'b0100000010100000000000000000000000000000011100000000000000000000;
mem[80] = 64'b0110010100100000000000000000000000000000000000000000000000000000;
mem[81] = 64'b0110010100100000000000000000000000000000000100000000000000000000;
mem[82] = 64'b0110010100100000000000000000000000000000001000000000000000000000;
mem[83] = 64'b0110010100100000000000000000000000000000001100000000000000000000;
mem[84] = 64'b0110010110000000000000000000000000000000010000000000000000000000;
mem[85] = 64'b0110010100100000000000000000000000000000010100000000000000000000;
mem[86] = 64'b0110010100100000000000000000000000000000011000000000000000000000;
mem[87] = 64'b0110010100100000000000000000000000000000011100000000000000000000;
mem[88] = 64'b0110000100000000000000000000000000000000010000000000000000000000;
mem[89] = 64'b0110000101100000000000000000000000000000010000000000000000000000;
mem[90] = 64'b0110000111000000000000000000000000000000010000000000000000000000;
mem[91] = 64'b0110001000100000000000000000000000000000010000000000000000000000;
mem[92] = 64'b0110001010000000000000000000000000000000010000000000000000000000;
mem[93] = 64'b0110001011100000000000000000000000000000010000000000000000000000;
mem[94] = 64'b0110001101000000000000000000000000000000010000000000000000000000;
mem[95] = 64'b0110001110100000000000000000000000000000010000000000000000000000;
mem[96] = 64'b0110011100100000000000000000000000000000010000000000000000000000;
mem[97] = 64'b0110100101000000000000000000000000000000010000000000000000000000;
mem[98] = 64'b0010110001100000000000000000000010010000000000000000110000000000;
mem[99] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[100] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[101] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[102] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[103] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[104] = 64'b0110011000100000000000000000000000000000010000000000000000000000;
mem[105] = 64'b0101101111100000000000000000000010010000100000000000110000000000;
mem[106] = 64'b0110011010000000000000000000000000000000010000000000000000000000;
mem[107] = 64'b0101101111100000000000000000000010010000100000000000110000000000;
mem[108] = 64'b0100100000000000000000000000000000000000000000000000000000000000;
mem[109] = 64'b0100100110100000000000000000000000000000000000000000000000000000;
mem[110] = 64'b0100010100000000000000000000000000000000000000000000000000000000;
mem[111] = 64'b0100011010000000000000000000000000000000000000000000000000000000;
mem[112] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[113] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[114] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[115] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[116] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[117] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[118] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[119] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[120] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[121] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[122] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[123] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[124] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[125] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[126] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[127] = 64'b0100110011100000000000000000000000000000000000000000000000000000;
mem[128] = 64'b1000011101100000000000000000000110010000000000000000000000000000;
mem[129] = 64'b1000011101100000000000000000000110010000000000000000000000000000;
mem[130] = 64'b1000011101100000000000000000000110010000000000000000000000000000;
mem[131] = 64'b1000100001100000000000000000000110010000000000000000000000000000;
mem[132] = 64'b1000000000100000000000000000000010010000100000000000110000000010;
mem[133] = 64'b1000000000100000000000000000000010010000100000000000110000000010;
mem[134] = 64'b1000000101100000000000000000000010010000100000000000110000000010;
mem[135] = 64'b1000000101100000000000000000000010010000100000000000110000000000;
mem[136] = 64'b0101001011100000000000000000000010010000000000000000000000000001;
mem[137] = 64'b0101001011100000000000000000000010010000000000000000000000000000;
mem[138] = 64'b0101001100100000000000000000000010010000100000000000110000000001;
mem[139] = 64'b0101001100100000000000000000000010010000100000000000110000000000;
mem[140] = 64'b0101010110000000000000000000000110010000000000000000000000000000;
mem[141] = 64'b0100111000000000000000000000000010010000000000000000110000000000;
mem[142] = 64'b0101010100100000000000000000000010010000100000000000110000000000;
mem[143] = 64'b1000100101100000000000000000000110010000000000000000100000000000;
mem[144] = 64'b0001001000100000000000000000000000000001000000000000000000000000;
mem[145] = 64'b1000001001000000000000000000000000000000000100000000000000000000;
mem[146] = 64'b1000001010100000000000000000000000000000001000000000000000000000;
mem[147] = 64'b1000001100000000000000000000000000000000001100000000000000000000;
mem[148] = 64'b1000001101100000000000000000000000000000010000000000000000000000;
mem[149] = 64'b1000001111000000000000000000000000000000010100000000000000000000;
mem[150] = 64'b1000010000100000000000000000000000000000011000000000000000000000;
mem[151] = 64'b1000010010000000000000000000000000000000011100000000000000000000;
mem[152] = 64'b0011110001100000000000000000000000000000000000000000000000000001;
mem[153] = 64'b0011110010000000000000000000000000000000000000000000000000000000;
mem[154] = 64'b0010111100000000001001000000000001001000000000000000010000000000;
mem[155] = 64'b0001001110000000000000000000000000000001000000000000000000000000;
mem[156] = 64'b0110011011100001011000000000000000001000010000000000000000000000;
mem[157] = 64'b0110010000000000000000000000000000000000010000000000000000000000;
mem[158] = 64'b0011110010100000000000000000000000000000010000000000000000000001;
mem[159] = 64'b0001010000000001011000000000000000000001000001001100000000000001;
mem[160] = 64'b0101010011000000001001000000000000110000000000000000110000000000;
mem[161] = 64'b0101010011000000001001000000000000110000000000000000110000000000;
mem[162] = 64'b0101010100000000001001000000000000110000000000000000000000000000;
mem[163] = 64'b0101010100000000001001000000000000110000000000000000000000000000;
mem[164] = 64'b0101011011000000000000000000000000000000000000000000000000000000;
mem[165] = 64'b0101100000100000000000000000000000000000000000000000000000000000;
mem[166] = 64'b0011001101100000000000000000000000000000000000000000000000000000;
mem[167] = 64'b0011010011100000000000000000000000000000000000000000000000000000;
mem[168] = 64'b1000000010000000000000000000000000000000000000000000000000000010;
mem[169] = 64'b1000000010000000000000000000000000000000000000000000000000000010;
mem[170] = 64'b0111101111100000000000000000000000000000000000000000000000000001;
mem[171] = 64'b0111110101000000000000000000000000000000000000000000000000000000;
mem[172] = 64'b0100111110000000000000000000000000000000000000000000000000000000;
mem[173] = 64'b0101000010000000000000000000000000000000000000000000000000000000;
mem[174] = 64'b0111011100100000000000000000000000000000011100000000000000000000;
mem[175] = 64'b0111100000100000000000000000000000000000011100000000000000000000;
mem[176] = 64'b0001011000100000001001000000000000000001000000001100000000000001;
mem[177] = 64'b0001011001000000001001000000000000000001000000011100000000000001;
mem[178] = 64'b0001011001100000001001000000000000000001000000101100000000000001;
mem[179] = 64'b0001011010000000001001000000000000000001000000111100000000000001;
mem[180] = 64'b0001011010100000001001000000000000000001000001001100000000000001;
mem[181] = 64'b0001011011000000001001000000000000000001000001011100000000000001;
mem[182] = 64'b0001011011100000001001000000000000000001000001101100000000000001;
mem[183] = 64'b0001011100000000001001000000000000000001000001111100000000000001;
mem[184] = 64'b0001011100100000001001000000000000000001000000001100000000000000;
mem[185] = 64'b0001011101000000001001000000000000000001000000011100000000000000;
mem[186] = 64'b0001011101100000001001000000000000000001000000101100000000000000;
mem[187] = 64'b0001011110000000001001000000000000000001000000111100000000000000;
mem[188] = 64'b0001011110100000001001000000000000000001000001001100000000000000;
mem[189] = 64'b0001011111000000001001000000000000000001000001011100000000000000;
mem[190] = 64'b0001011111100000001001000000000000000001000001101100000000000000;
mem[191] = 64'b0001100000000000001001000000000000000001000001111100000000000000;
mem[192] = 64'b1000101101100000000000000000000110010000000000000000000000000001;
mem[193] = 64'b1000110001100000000000000000000110010000000000000000000000000000;
mem[194] = 64'b0110111001000000000000000000000000000000010000000000000000000000;
mem[195] = 64'b0110110111100000000000000000000000000000010000000000000000000000;
mem[196] = 64'b0100111011000000000000000000000010010000000000000000110000000000;
mem[197] = 64'b0100110101000000000000000000000010010000000000000000110000000000;
mem[198] = 64'b0101001110000000000000000000000110010000000000000000000000000000;
mem[199] = 64'b0101001110000000000000000000000110010000000000000000000000000000;
mem[200] = 64'b0011100111100000001001000000000000000000010000000000000010000000;
mem[201] = 64'b0100111001000000000000000000000000000000010100000000000000000000;
mem[202] = 64'b0110111101100000000000000000000000000000010000000000000000000000;
mem[203] = 64'b0110111011000000000000000000000000000000010000000000000000000000;
mem[204] = 64'b0010010110100000001001000111000000000000000000000000000010000000;
mem[205] = 64'b0100000011000000001001000000000000110000000000000000000000000000;
mem[206] = 64'b0100000100000001011000000000000000001000000000000000000000000000;
mem[207] = 64'b0111000000100000000000000000000000000000010000000000000000000000;
mem[208] = 64'b1000101001100000000000000000000110010000000000000000000000000010;
mem[209] = 64'b1000101001100000000000000000000110010000000000000000000000000000;
mem[210] = 64'b1000110101100000000000000000000110010000000000000000000000000010;
mem[211] = 64'b1000110101100000000000000000000110010000000000000000000000000000;
mem[212] = 64'b0011100100000000001001000000000000001000100000000000000000000001;
mem[213] = 64'b0010011000100000000000000000000000000000010000000000000000000001;
mem[214] = 64'b0011110011000000000000000000000000000000000110000000000000000000;
mem[215] = 64'b1000010011100000000000000000000000000000000000000000000000000001;
mem[216] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[217] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[218] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[219] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[220] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[221] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[222] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[223] = 64'b0011110001000000000000000000000000000000000000000000000000000000;
mem[224] = 64'b0101001010000000000000000000000000000000000100000000000000000000;
mem[225] = 64'b0101001000000000000000000000000000000000000100000000000000000000;
mem[226] = 64'b0101000110000000000000000000000000000000000100000000000000000000;
mem[227] = 64'b0100110010000000000000000000000000000000000010000000000000000000;
mem[228] = 64'b0100010001000000001001000000000000110000000000000000000000000001;
mem[229] = 64'b0100010001000000001001000000000000110000000000000000000000000001;
mem[230] = 64'b0100001110000000001001000000000000110000000000000000000000000001;
mem[231] = 64'b0100001110000000001001000000000000110000000000000000000000000001;
mem[232] = 64'b0010110111100000000000000000000000000000010000000000000000000000;
mem[233] = 64'b0001110101001000010001000000000001000001000000000000000000000000;
mem[234] = 64'b0100101101000000001001000000000001000000000000000000000000000000;
mem[235] = 64'b0001110110001000010001000000000001000001000000000000000000000000;
mem[236] = 64'b0100010010100000000000000000000000000000001000000000000000000000;
mem[237] = 64'b0100010010100000000000000000000000000000001000000000000000000000;
mem[238] = 64'b0100001111100000000000000000000000000000000000000000000000000001;
mem[239] = 64'b0100001111100000000000000000000000000000000000000000000000000000;
mem[240] = 64'b0001111000100000000000000000000000000001000000000000000000000000;
mem[241] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[242] = 64'b0001111001100000000000000000000000000001000000000000000000000000;
mem[243] = 64'b0001111010000000000000000000000000000001000000000000000000000000;
mem[244] = 64'b0011110011100000000000000000000000000000000000000000000000000000;
mem[245] = 64'b0001111011000001110000000000000000000001000000000000000000010100;
mem[246] = 64'b1000111001100000000000000000000110010000000000000000000000000001;
mem[247] = 64'b1000111101100000000000000000000110010000000000000000000000000000;
mem[248] = 64'b0001111100100001100001000001000000000001000000000000000000010100;
mem[249] = 64'b0001111101000001100001000110000000000001000000000000000000010100;
mem[250] = 64'b0001111101100001100001100001000000000001000000000000000000011100;
mem[251] = 64'b0001111110000001100001100110000000000001000000000000000000011100;
mem[252] = 64'b0001111110100001100001000001000000000001000000000000000000100000;
mem[253] = 64'b0001111111000001100001000110000000000001000000000000000000100000;
mem[254] = 64'b0011110100000000000000000000000110010000000000000000000000000001;
mem[255] = 64'b1001000001100000000000000000000110010000000000000000110000000000;
mem[256] = 64'b0010000000100000000000010000000100000000000000000000000000000000;
mem[257] = 64'b0010010110100000001001000001000000000000000000000000000010000000;
mem[258] = 64'b0010000001000000000000000000000000000000000000000000000000000000;
mem[259] = 64'b1001001101000000000000000000000000000000000000000000000000000000;
mem[260] = 64'b1001001101000000000000000000000000000000000100000000000000000000;
mem[261] = 64'b1001001101000000000000000000000000000000001000000000000000000000;
mem[262] = 64'b1001001101000000000000000000000000000000001100000000000000000000;
mem[263] = 64'b1001001101000000000000000000000000000000010000000000000000000000;
mem[264] = 64'b1001001101000000000000000000000000000000010100000000000000000000;
mem[265] = 64'b1001001101000000000000000000000000000000011000000000000000000000;
mem[266] = 64'b1001001101000000000000000000000000000000011100000000000000000000;
mem[267] = 64'b1001001101100000000000000000000000000000000000000000001000000000;
mem[268] = 64'b1001001101100000000000000000000000000000000000000000011000000000;
mem[269] = 64'b1001001101100000000000000000000000000000000000000000101000000000;
mem[270] = 64'b1001001101100000000000000000000000000000000000000000111000000000;
mem[271] = 64'b0010000001001000000000000000000000000000000000000000000010000000;
mem[272] = 64'b0010000001000001011000000000000000000000000000000000000010000000;
mem[273] = 64'b0010000001000000001011100000000001000001000000000000000000000000;
mem[274] = 64'b0010000001000001100011000000000000000000000000000000000000110000;
mem[275] = 64'b0010000001000000001011000000000000000000000000001100000000000000;
mem[276] = 64'b0010000001000000001011000000000000000000000000011100000000000000;
mem[277] = 64'b0010000001000000001011000000000000000000000000101100000000000000;
mem[278] = 64'b0010000001000000001011000000000000000000000000111100000000000000;
mem[279] = 64'b0010000001000000001011000000000000000000000001001100000000000000;
mem[280] = 64'b0010000001000000001011000000000000000000000001011100000000000000;
mem[281] = 64'b0010000001000000001011000000000000000000000001101100000000000000;
mem[282] = 64'b0010000001000000001011000000000000000000000001111100000000000000;
mem[283] = 64'b0010000001000000001011100000000000000001000000000000001100000000;
mem[284] = 64'b0010000001000000001011100000000000000001000000000000011100000000;
mem[285] = 64'b0010000001000000001011100000000000000001000000000000101100000000;
mem[286] = 64'b0010000001000000001011100000000000000001000000000000111100000000;
mem[287] = 64'b0010000001000000001011000000000000110000000000000000000000000000;
mem[288] = 64'b0010000001000000001011000000000000001000000000000000000000000000;
mem[289] = 64'b1001001110000000000000000000000000000000000000000000111000000000;
mem[290] = 64'b1001001111100000000000000000000000000000000000000000111000000000;
mem[291] = 64'b1001010001000000000000000000000000000000000000000000111000000000;
mem[292] = 64'b1001010010000000000000000000000000000000000000000000111000000000;
mem[293] = 64'b1001010011000000000000000000000000000000000000000000111000000000;
mem[294] = 64'b1001010100000000000000000000000000000000000000000000111000000000;
mem[295] = 64'b1001010101000000000000000000000000000000000000000000111000000000;
mem[296] = 64'b1001010101100000000000000000000000000000000000000000111000000000;
mem[297] = 64'b1001000101100000000000000000000000000000000000000000000000000000;
mem[298] = 64'b0010010110100000001001001011000000000000000000000000000010000000;
mem[299] = 64'b0010010110111011100001001001000000000000000000000000000010000000;
mem[300] = 64'b0010010110100000001001001001000000000000000000000000000010000000;
mem[301] = 64'b0100000101100001011000000000000000001000010000000000000000000000;
mem[302] = 64'b0010010111100000000000000000000100000000000000000000000000000000;
mem[303] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[304] = 64'b0010011000100011000000000000000000000001000000001100000000000100;
mem[305] = 64'b0010011001000011101001000000000000000000000000000000000010000000;
mem[306] = 64'b0010011001100000000000000000000000000000000000000000000000000001;
mem[307] = 64'b0010011010000000010011000000000000000000000000001100000000001000;
mem[308] = 64'b0010011010100000001001000001000000000001000001001100000000000001;
mem[309] = 64'b0010011011000011001000000000000000000001000000001100000000000100;
mem[310] = 64'b0010011011100000011000000000000000000001000000001000000000001110;
mem[311] = 64'b0010011100000000000000000000000000000100000000000000110000000010;
mem[312] = 64'b1001001100111000011000000000000000001000000000000000110000001110;
mem[313] = 64'b0010011101000000011000000000000000000001000000000100000000001110;
mem[314] = 64'b0010011101100000000000000000000000000100000000000000110000000010;
mem[315] = 64'b0010011110011000011000000000000000000001000000000100000000001110;
mem[316] = 64'b0010011110100000011001000000000000000001000000001100000000001110;
mem[317] = 64'b0010011111000000011001000000000000000001000000001000000000001110;
mem[318] = 64'b0010011111100000000000000000000000000100000000000000110000000010;
mem[319] = 64'b1001001100111000011001000000000000001000000000000000110000001110;
mem[320] = 64'b0010100001000000000000000000000000000000100000000000000000000000;
mem[321] = 64'b0010100001100000000000000000000000000000100000000000110000000000;
mem[322] = 64'b0010100001100000011001000000000000000001000000001000000000001100;
mem[323] = 64'b0010100010000000000000000000000000000100000000000000110000000000;
mem[324] = 64'b1001001100011000011001000000000000001000000000000000110000001100;
mem[325] = 64'b0010100011000000010000000000000000000001000000001000000000001110;
mem[326] = 64'b0010100011100000000000000000000000000100000000000000110000000010;
mem[327] = 64'b1001001100111000010000000000000000001000000000000000110000001110;
mem[328] = 64'b0010100100100000010000000000000000000001000000000100000000001110;
mem[329] = 64'b0010100101000000000000000000000000000100000000000000110000000010;
mem[330] = 64'b0010100101111000010000000000000000000001000000000100000000001110;
mem[331] = 64'b0010100110000000010001000000000000000001000000001100000000001110;
mem[332] = 64'b0010100110100000010001000000000000000001000000001000000000001110;
mem[333] = 64'b0010100111000000000000000000000000000100000000000000110000000010;
mem[334] = 64'b1001001100111000010001000000000000001000000000000000110000001110;
mem[335] = 64'b0010101000100000000000000000000000000000100000000000000000000000;
mem[336] = 64'b0010101001000000000000000000000000000000100000000000110000000000;
mem[337] = 64'b0010101001000000010001000000000000000001000000001000000000001100;
mem[338] = 64'b0010101001100000000000000000000000000100000000000000110000000000;
mem[339] = 64'b1001001100011000010001000000000000001000000000000000110000001100;
mem[340] = 64'b0010101010100000100000000000000000000001000000001000000000010010;
mem[341] = 64'b0010101011000000000000000000000000000100000000000000110000000010;
mem[342] = 64'b1001001100111000100000000000000000001000000000000000110000010010;
mem[343] = 64'b0010101100000000100000000000000000000001000000000100000000010010;
mem[344] = 64'b0010101100100000000000000000000000000100000000000000110000000010;
mem[345] = 64'b0010101101011000100000000000000000000001000000000100000000010010;
mem[346] = 64'b0010101101100000100001000000000000000001000000001100000000010010;
mem[347] = 64'b0010101110000000100001000000000000000001000000001000000000010010;
mem[348] = 64'b0010101110100000000000000000000000000100000000000000110000000010;
mem[349] = 64'b1001001100111000100001000000000000001000000000000000110000010010;
mem[350] = 64'b0010110000000000000000000000000000000000100000000000000000000000;
mem[351] = 64'b0010110000100000000000000000000000000000100000000000110000000000;
mem[352] = 64'b0010110000100000100001000000000000000001000000001000000000010000;
mem[353] = 64'b0010110001000000000000000000000000000100000000000000110000000000;
mem[354] = 64'b1001001100011000100001000000000000001000000000000000110000010000;
mem[355] = 64'b0010010110100000001001000010000000000000000000000000000010000000;
mem[356] = 64'b0010110010100001011000000000000000000100000000000000110010000000;
mem[357] = 64'b0010110011011100001000000000000000000000000000000000000000010100;
mem[358] = 64'b0010110101110000010001000011001110110000000000000000110000000000;
mem[359] = 64'b0010110100000000000000000000000000000100000000000000110000000000;
mem[360] = 64'b0010110100111100010000000000000000000000000000000000000000010100;
mem[361] = 64'b0010110101100000000000000000001110000000000000000000000000000000;
mem[362] = 64'b0010110101100001100011000000000000000001000000000000000000010100;
mem[363] = 64'b0010110110000001100011000000000000000000000000000000000000010100;
mem[364] = 64'b0010010110100000001001000100000000000000000000000000000010000000;
mem[365] = 64'b0010110111000011010000000000000000000001000000001100000000011000;
mem[366] = 64'b0010110111100011011000000000000000000001000000001100000000011000;
mem[367] = 64'b0010111000000000111001000011000000110000000001001100000000000000;
mem[368] = 64'b0010111000101000000000000000000000001000010000000000101000000000;
mem[369] = 64'b0010111001001000010001000000000001000011000000000000101000000000;
mem[370] = 64'b0010111010100000000000000000000001000000010000000000000000000000;
mem[371] = 64'b0010111010000000000000000000000000000100000000000000110000000000;
mem[372] = 64'b0010111010111000000000000000000001000000010000000000000000000000;
mem[373] = 64'b0010111011000000111001000011000000110000000001001100000000000000;
mem[374] = 64'b0010111011101000000000000000000000001000010000000000101000000000;
mem[375] = 64'b0010111100000000000000000000000000000011000000000000101000000000;
mem[376] = 64'b0010111100100000001010000000000000001000010000000000000000000000;
mem[377] = 64'b0010111101000000111001000011000000110000000001001100101000000000;
mem[378] = 64'b0010111101100000000000000000000000000010010000000000101000000000;
mem[379] = 64'b0010111110000000111001000011000000110000000001001100000000000000;
mem[380] = 64'b0010111110101000000000000000000000001000000000000000101000000000;
mem[381] = 64'b0010111111000000000000000000000000000010000000000000101000000000;
mem[382] = 64'b0010111111100000001100000000000000000001000000000000011100000000;
mem[383] = 64'b0011000000000000000000000000000000000001000000000000000000000000;
mem[384] = 64'b0011000000100000001010000000000000001000010000000000000000000000;
mem[385] = 64'b0011000001000000111001000011000000110000000001001100101000000000;
mem[386] = 64'b0011000001100000000000000000000000000010010000000000101000000000;
mem[387] = 64'b0011000010000000111001000011000000110000000001001100000000000000;
mem[388] = 64'b0011000010101000000000000000000000001000000000000000101000000000;
mem[389] = 64'b0011000011000000000000000000000000000010000000000000101000000000;
mem[390] = 64'b0011000011100000000000000000000000010000000000000000110000000000;
mem[391] = 64'b0011000100000000000000000000000000000100000000000000110000000000;
mem[392] = 64'b0011000100111000000000000000000001000000000000000000000000000000;
mem[393] = 64'b0011000101010000010001000011000000110000000000000000110000000000;
mem[394] = 64'b0011000101100000000000000000000000000100000000000000110000000000;
mem[395] = 64'b0011000110011000000000000000000000000001000000000000011100000000;
mem[396] = 64'b0011000110100000111000000000000000000001000000000000000000001110;
mem[397] = 64'b0011000111000000000000000000000000000100000000000000110000000010;
mem[398] = 64'b0011000111111000111000000000000000000001000000000000000000001110;
mem[399] = 64'b0011001000000001000000000000000000000001000000000000000000001110;
mem[400] = 64'b0011001000100000000000000000000000000100000000000000110000000010;
mem[401] = 64'b0011001001011001000000000000000000000001000000000000000000001110;
mem[402] = 64'b0011001001100000111001000000000000000001000000000000000000001110;
mem[403] = 64'b0011001010000000111001000000000000000001000000000000000000001110;
mem[404] = 64'b0011001010100000000000000000000000000100000000000000110000000010;
mem[405] = 64'b0011001011011000111001000000000000000001000000000000000000001110;
mem[406] = 64'b0011001100000000000000000000000000000000100000000000000000000000;
mem[407] = 64'b0011001100100000000000000000000000000000100000000000110000000000;
mem[408] = 64'b0011001100100000111001000000000000000001000000000000000000001100;
mem[409] = 64'b0011001101000000000000000000000000000100000000000000110000000000;
mem[410] = 64'b0011001101111000111001000000000000000001000000000000000000001100;
mem[411] = 64'b0011001111000000000000000000001000000000011110000000000000000000;
mem[412] = 64'b0011010011000000000000000000010000000000000100000000000000000000;
mem[413] = 64'b0011001111000000111001000101000000000000011100011100000000000000;
mem[414] = 64'b0011001111100000000000000000000000110000011100000000001000000000;
mem[415] = 64'b0011010000011000000000000000000000000100000000000000001010000001;
mem[416] = 64'b0011010000110010111001000101000000000000011001111100000000000000;
mem[417] = 64'b0011010001000000000000000000000000110000011000000000110000000000;
mem[418] = 64'b0011010001100010111001000101000000000000000001101100110000000000;
mem[419] = 64'b0011010010000000000000000000000000000100000000000000110000000001;
mem[420] = 64'b0011010011011000111011000000001000000000000000000000000000001101;
mem[421] = 64'b0011001110000001011000010000001100000000000010000000000000000000;
mem[422] = 64'b0011010011100000000000000000000000000001000000000000000000000000;
mem[423] = 64'b0011010101000000000000000000001000000000011110000000000000000000;
mem[424] = 64'b0011011000100000000000000000010000000000000100000000000000000000;
mem[425] = 64'b0011010101000000111001000101000000000000011100011100000000000000;
mem[426] = 64'b0011010101100000000000000000000000110000011100000000001000000000;
mem[427] = 64'b0011010110011000000000000000000000000100011100000000001010000000;
mem[428] = 64'b0011010110100010111001000011000000000000011001111100000000000000;
mem[429] = 64'b0011010111000000000000000000000000110000011000000000110000000000;
mem[430] = 64'b0011010111100010111001000011000000000000000001101100110000000000;
mem[431] = 64'b0011011000111000111011000000001000000100000000000000110000001100;
mem[432] = 64'b0011010100000001011000010000001100000000000010000000000000000000;
mem[433] = 64'b0011011001000000000000000000000000000001000000000000000000000000;
mem[434] = 64'b0011011010000000000000000000000000001000000000000000000000000001;
mem[435] = 64'b0011011010000000000000000000000000000100000000000000110000000001;
mem[436] = 64'b0011011010100000000000000000000000000000000000000000000000000000;
mem[437] = 64'b0011011011000000000000000000000000000000000000000000000010000000;
mem[438] = 64'b0011011011100011110000000000000000000000000000000000000000000001;
mem[439] = 64'b0011011100000000000000000000000000000000000000001101000000000001;
mem[440] = 64'b0011011100100000000000000000000000000001000001001110000000000001;
mem[441] = 64'b0011011101100000000000000000000000001000000000000000000000000000;
mem[442] = 64'b0011011101100000000000000000000000000100000000000000110000000000;
mem[443] = 64'b0011011110000000000000000000000000000000001000000000000010000000;
mem[444] = 64'b0011011110100011110000000000000000000000001000000000000000000000;
mem[445] = 64'b0011011111000000000000000000000000000000000000001101000000000000;
mem[446] = 64'b0011011111100000000000000000000000000001000000101110000000000000;
mem[447] = 64'b0011100000100000000000000000000000001000000000000000000000000001;
mem[448] = 64'b0011100000100000000000000000000000000100000000000000110000000001;
mem[449] = 64'b0011100001000000000000000000000000000000000000000000000000000000;
mem[450] = 64'b0011100001100000000000000000000000000000000000000000000010000000;
mem[451] = 64'b0011011011100011111000000000000000000000000000000000000000000001;
mem[452] = 64'b0011100011000000000000000000000000001000000000000000000000000000;
mem[453] = 64'b0011100011000000000000000000000000000100000000000000110000000000;
mem[454] = 64'b0011100011100000000000000000000000000000001000000000000010000000;
mem[455] = 64'b0011011110100011111000000000000000000000001000000000000000000000;
mem[456] = 64'b0011100100100000000000000000000000000000000000000000000000000001;
mem[457] = 64'b0011100101000000000000000000000000000000000000000000000010000000;
mem[458] = 64'b0011100101100011110000000000000000000000000000000000000000000001;
mem[459] = 64'b0011100110000000000000000000000000000000000001001101000000000001;
mem[460] = 64'b0011100110100000000000000000000000000000000000001110000000000001;
mem[461] = 64'b0011100111000000000000000000000000000000000000000000000000000000;
mem[462] = 64'b0011100111100000010001000001000000000001000000000000000000001000;
mem[463] = 64'b0011101000000000111001000011000000110000010101001100000000000000;
mem[464] = 64'b0011101000100000000000000000000000001000000000000000101000000000;
mem[465] = 64'b0011110000000000000000000000010010000010010000000000101000000000;
mem[466] = 64'b0011101001100100011100000000000000110000010000000000000000000000;
mem[467] = 64'b0011101010000000000000000000000000001000000000000000101000000000;
mem[468] = 64'b0011101010100000000000000000000000000010000000000000101000000000;
mem[469] = 64'b0011101101100000000000000000010010000000010100000000000000000000;
mem[470] = 64'b0011101011100000111001000011000000110000000001011100101000000000;
mem[471] = 64'b0011101100000000000000000000000000000100010000000000101000000000;
mem[472] = 64'b0011101100100000111001000011000000110000000001001100101000000000;
mem[473] = 64'b0011101101000000000000000000000000000010000000000000101000000000;
mem[474] = 64'b0011101010100000000000000000000000000000000000000000000000000000;
mem[475] = 64'b0011101110000000000000000000000000000000010000000000000000000000;
mem[476] = 64'b0011101110100000111001000011000000110000000001001100101000000000;
mem[477] = 64'b0011101111000000000000000000000000000100010000000000101000000000;
mem[478] = 64'b0011101111111000000000000000000000000000010001011100000000000000;
mem[479] = 64'b0011110000000000111011000000000000000001000001001100000000000000;
mem[480] = 64'b0011110000100000000000000000000000000000010001011100000000000000;
mem[481] = 64'b0011110001000000111011000000000000000001000001001100000000000000;
mem[482] = 64'b0011110001100000000000000000000000000001000000000000000000000000;
mem[483] = 64'b0011110010000100000001000000000000000001000001001100000000000001;
mem[484] = 64'b0011110010100100000001000000000000000001000000101100000000000000;
mem[485] = 64'b0011110011000001101000000000000000000001000000000000000000011000;
mem[486] = 64'b0011110011100001001000000000000000000001000000001100000000000001;
mem[487] = 64'b0011110011100000000000010000000000000000000000000000000000000000;
mem[488] = 64'b0011111000000000000000000000000010000000100000000000110000000001;
mem[489] = 64'b0011111001100000000000000000000010000000100000000000110000000001;
mem[490] = 64'b0011110101100000000000000000000000000001000000000000000000000000;
mem[491] = 64'b0011110110000000000000000000000000000001000000000000000000000000;
mem[492] = 64'b0011110110100000000000000000000000000001000000000000000000000000;
mem[493] = 64'b0011110111000000000000000000000000000001000000000000000000000000;
mem[494] = 64'b0011110111100000000000000000000000000001000000000000000000000000;
mem[495] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[496] = 64'b0011111000100000010001000101000000000001000000001000000000100110;
mem[497] = 64'b0011111001000000000000000000000000000100000000000000110000000010;
mem[498] = 64'b1001001100111000010001000101000000001000000000000000110000100110;
mem[499] = 64'b0011111010000000111001000101000000000001000000001000000000100110;
mem[500] = 64'b0011111010100000000000000000000000000100000000000000110000000010;
mem[501] = 64'b1001001100111000111001000101000000001000000000000000110000100110;
mem[502] = 64'b0011111011100000010001000101000000000001000000001100000000100100;
mem[503] = 64'b0011111100000000010001000101000000000001000000011100000000100100;
mem[504] = 64'b0011111100100000010001000101000000000001000000101100000000100100;
mem[505] = 64'b0011111101000000010001000101000000000001000000111100000000100100;
mem[506] = 64'b0011111101100000010001000101000000000001000001001100000000100100;
mem[507] = 64'b0011111110000000010001000101000000000001000001011100000000100100;
mem[508] = 64'b0011111110100000010001000101000000000001000001101100000000100100;
mem[509] = 64'b0011111111000000010001000101000000000001000001111100000000100100;
mem[510] = 64'b0011111111100000111001000101000000000001000000001100000000100100;
mem[511] = 64'b0100000000000000111001000101000000000001000000011100000000100100;
mem[512] = 64'b0100000000100000111001000101000000000001000000101100000000100100;
mem[513] = 64'b0100000001000000111001000101000000000001000000111100000000100100;
mem[514] = 64'b0100000001100000111001000101000000000001000001001100000000100100;
mem[515] = 64'b0100000010000000111001000101000000000001000001011100000000100100;
mem[516] = 64'b0100000010100000111001000101000000000001000001101100000000100100;
mem[517] = 64'b0100000011000000111001000101000000000001000001111100000000100100;
mem[518] = 64'b0100000011110000100001001000000000110000000000000000000000000000;
mem[519] = 64'b0010010110110011100001001001000000000000000000000000000010000000;
mem[520] = 64'b0100000101000000001001001010001110000000010000000000000010000000;
mem[521] = 64'b0100000101000000000000000000000000000001000000000000000000000000;
mem[522] = 64'b0010010110100000000000000000000000000000000000000000000000000000;
mem[523] = 64'b0100000110000000111001000011000000110000000000000000101000000000;
mem[524] = 64'b0100000110100000000000000000000000000010000000000000101000000000;
mem[525] = 64'b0100000111010000111001000011000000110000000000000000011000000000;
mem[526] = 64'b0100000111100000001010000000000000001000000000000000101000000000;
mem[527] = 64'b0100001000000000000000000000000000000010000000000000101000000000;
mem[528] = 64'b0100001000110000111001000011000000110000000000000000000000000000;
mem[529] = 64'b0100001001001000000000000000000000001000000000000000101000000000;
mem[530] = 64'b0100001001100000000000000000000000000010000000000000101000000000;
mem[531] = 64'b0100001010010000000000000000000000000000000001001100000000000000;
mem[532] = 64'b0100001010100001100001000001000000000000000000000000000000101000;
mem[533] = 64'b0100001011000000001001000001000000000000000000000000011100000000;
mem[534] = 64'b0100001011100000001011000000000000110000000000000000011000000000;
mem[535] = 64'b0100001100000000000000000000000000000100000000000000011000000000;
mem[536] = 64'b0100001100111000000000000000000001000000000000000000000000000000;
mem[537] = 64'b0100001101010000010001000011000000110000000000000000011000000000;
mem[538] = 64'b0100001101100000000000000000000000000100000000000000011000000000;
mem[539] = 64'b0100001110011000000000000000000000000001000000000000011100000000;
mem[540] = 64'b0100001110110000100001001000000000110000000000000000000000000000;
mem[541] = 64'b0100001111000000000000000000000000001000000000000000000000000000;
mem[542] = 64'b0100001111100000000000000000100000000011000000000000000000000010;
mem[543] = 64'b0100010000000000000000000000000000001000001000000000000000000000;
mem[544] = 64'b0100010000100000000000000000000000110000000000000000000000000000;
mem[545] = 64'b0100010001000000000000000000100000000011000000000000000000000010;
mem[546] = 64'b0100010001110000100001001000000000110000000000000000000000000000;
mem[547] = 64'b0100010010000000000000000000100000000100000000000000000000000010;
mem[548] = 64'b0100010010111000000000000000000000000001000000001100000000000010;
mem[549] = 64'b0100010011000000000000000000000000110000000000000000000000000000;
mem[550] = 64'b0100010011100000000000000000100000000100000000000000000000000010;
mem[551] = 64'b0100010100011000000000000000000000000001000000001100000000000010;
mem[552] = 64'b0100010110000000000000000000001000000000011000000000000000000000;
mem[553] = 64'b0100010101000000000000000000000000000000000010000000000000000000;
mem[554] = 64'b0100011001100000111001000001010000000000000100000000000000000000;
mem[555] = 64'b0100010110000000111001000101000000000000011000011100000000000000;
mem[556] = 64'b0100010110100000000000000000000000110000011000000000110000000000;
mem[557] = 64'b0100010111000010111001000101000000000000000001101100110000000000;
mem[558] = 64'b0100010111100000000000000000000000000100000000000000110000000001;
mem[559] = 64'b0100011000000000000000000000000000000000001000000000000000000000;
mem[560] = 64'b0100011000100000000000000000000000110000000000000000000000000000;
mem[561] = 64'b0100011001100000000000000000101000000010000000000000000000000001;
mem[562] = 64'b0100010101000000000000010000000000000000000010000000000000000000;
mem[563] = 64'b0100011010000000000000000000000000000001000000000000000000000000;
mem[564] = 64'b0100011100000000000000000000001000000000011000000000000000000000;
mem[565] = 64'b0100011011000000000000000000000000000000000010000000000000000000;
mem[566] = 64'b0100011111100000111001000001010000000000000100000000000000000000;
mem[567] = 64'b0100011100000000111001000101000000000000011000011100000000000000;
mem[568] = 64'b0100011100100000000000000000000000110000011000000000110000000000;
mem[569] = 64'b0100011101000010111001000011000000000000000001101100110000000000;
mem[570] = 64'b0100011101100000000000000000000000000100000000000000110000000000;
mem[571] = 64'b0100011110000000000000000000000000000000001000000000000000000000;
mem[572] = 64'b0100011110100000000000000000000000110000000000000000000000000000;
mem[573] = 64'b0100011111100000000000000000101000000010000000000000000000000000;
mem[574] = 64'b0100011011000000000000010000000000000000000010000000000000000000;
mem[575] = 64'b0100100000000000000000000000000000000001000000000000000000000000;
mem[576] = 64'b0100100010000000000000000000001000000000001000000000000000000000;
mem[577] = 64'b0100100001000000000000000000000000000000000010000000000000000000;
mem[578] = 64'b0100100110000000111001000001010000000000000100000000000000000000;
mem[579] = 64'b0100100010000000111001000101000000000000001000011100000000000000;
mem[580] = 64'b0100100010100000000000000000000000110000000000000000000000000000;
mem[581] = 64'b0100100011000000000000000000100000000100000000000000000000000001;
mem[582] = 64'b0100100011100000000000000000000000000000011100000000000000000000;
mem[583] = 64'b0100100100000000000000000000000000110000000000000000001000000000;
mem[584] = 64'b0100100100100000000000000000000000000010000000000000001000000001;
mem[585] = 64'b0100100101000000000000000000000000000000011100000000000000000000;
mem[586] = 64'b0100100110000010111001000101001000000000000001111100000000000000;
mem[587] = 64'b0100100001000000000000010000000000000000000010000000000000000000;
mem[588] = 64'b0100100110100000000000000000000000000001000000000000000000000000;
mem[589] = 64'b0100101000100000000000000000001000000000001000000000000000000000;
mem[590] = 64'b0100100111100000000000000000000000000000000010000000000000000000;
mem[591] = 64'b0100101100100000111001000001010000000000000100000000000000000000;
mem[592] = 64'b0100101000100000111001000101000000000000001000011100000000000000;
mem[593] = 64'b0100101001000000000000000000000000110000000000000000000000000000;
mem[594] = 64'b0100101001100000000000000000100000000100000000000000000000000000;
mem[595] = 64'b0100101010000000000000000000000000000000011100000000000000000000;
mem[596] = 64'b0100101010100000000000000000000000110000000000000000001000000000;
mem[597] = 64'b0100101011000000000000000000000000000010000000000000001000000000;
mem[598] = 64'b0100101011100000000000000000000000000000011100000000000000000000;
mem[599] = 64'b0100101100100010111001000011001000000000000001111100000000000000;
mem[600] = 64'b0100100111100000000000010000000000000000000010000000000000000000;
mem[601] = 64'b0100101101000000000000000000000000000001000000000000000000000000;
mem[602] = 64'b0100101101100000001100000000000000000001000000000000011100000000;
mem[603] = 64'b0100101110000000000000000000000001000001000000000000000000000000;
mem[604] = 64'b0100101110100000000000000000000000000100000000000000110000000000;
mem[605] = 64'b0100101111011000000000000000000001000001000000000000000000000000;
mem[606] = 64'b0100101111100000000000000000000000000001000000000000000000000000;
mem[607] = 64'b0100110000000000000000000000000000000100000000000000110000000000;
mem[608] = 64'b0100110000111000000000000000000001000000000000000000000000000000;
mem[609] = 64'b0100110001010000010001000011000000110000000000000000110000000000;
mem[610] = 64'b0100110001100000000000000000000000000100000000000000110000000000;
mem[611] = 64'b0100110010011000000000000000000000000001000000000000011100000000;
mem[612] = 64'b0100110011000000000000000000010000000000000000000000000000000000;
mem[613] = 64'b0100110011000000000000000000000000000001000000000000000000000000;
mem[614] = 64'b0100110011101000010001000000000001000001000000000000000000000000;
mem[615] = 64'b0100110100100000000000000000001110000000000000000000000000000000;
mem[616] = 64'b0100110100100000000000000000000000000001000000000000000000000000;
mem[617] = 64'b0100110101001000010001000000000001000001000000000000000000000000;
mem[618] = 64'b0100110101100000000000000000000000000001000000000000000000000000;
mem[619] = 64'b0100110110000000000000000000000000000100000000000000110000000000;
mem[620] = 64'b0100110110111000000000000000000000000000000000000100110000000000;
mem[621] = 64'b0100110111010000010001000011000000110000000000000000110000000000;
mem[622] = 64'b0100110111100000000000000000000000000100000000000000110000000000;
mem[623] = 64'b0100111000011000000000000000000000000001000000000000111100000000;
mem[624] = 64'b0100111000100000000000000000000000000001000000000000000000000000;
mem[625] = 64'b0100111001010000000000000000000000000001000000000100000000000000;
mem[626] = 64'b0100111001100000000000000000000000110000000001001100101000000000;
mem[627] = 64'b0100111010000000000000000000000000000100000000000000101000000000;
mem[628] = 64'b0100111010111000000000000000000000000000000001011100000000000000;
mem[629] = 64'b0100111011010000010001000011000000000001000001001100000000000000;
mem[630] = 64'b0100111011100000000000000000000000000001000000000000000000000000;
mem[631] = 64'b0100111100000000000000000000000000000100000000000000110000000000;
mem[632] = 64'b0100111100111000000000000000000000000000000000000100110000000000;
mem[633] = 64'b0100111101010000010001000011000000110000000000000000110000000000;
mem[634] = 64'b0100111101100000000000000000000000000100000000000000110000000000;
mem[635] = 64'b0100111110011000000000000000000000000001000000000000001100000000;
mem[636] = 64'b0100111111100000000000000000001000000000011010000000000000000000;
mem[637] = 64'b0101000001100000000000000000010000000000000100000000000000000000;
mem[638] = 64'b0100111111100000111001000101000000000000011000011100000000000000;
mem[639] = 64'b0101000000000000000000000000000000110000011000000000110000000000;
mem[640] = 64'b0101000000100010111001000101000000000000000001101100110000000000;
mem[641] = 64'b0101000001111000000000000000001000000100000000001100110000000001;
mem[642] = 64'b0100111110100000000000010000000000000000000010000000000000000000;
mem[643] = 64'b0101000010000000000000000000000000000001000000000000000000000000;
mem[644] = 64'b0101000011100000000000000000001000000000011010000000000000000000;
mem[645] = 64'b0101000101100000000000000000010000000000000100000000000000000000;
mem[646] = 64'b0101000011100000111001000101000000000000011000011100000000000000;
mem[647] = 64'b0101000100000000000000000000000000110000011000000000110000000000;
mem[648] = 64'b0101000100100010111001000011000000000000000001101100110000000000;
mem[649] = 64'b0101000101111000000000000000001000000100000000001100110000000000;
mem[650] = 64'b0101000010100000000000010000000000000000000010000000000000000000;
mem[651] = 64'b0101000110000000000000000000000000000001000000000000000000000000;
mem[652] = 64'b0101000110100000111001000101000000000000000010011100000000000000;
mem[653] = 64'b0101000111100000000000000000010000000000000000000000000000000000;
mem[654] = 64'b0101000111101000010001000000000001000001000000000000000000000000;
mem[655] = 64'b0101001000000000000000000000000000000001000000000000000000000000;
mem[656] = 64'b0101001001000000111001000101001010000000000010011100000000000000;
mem[657] = 64'b0101000111100000000000000000000000000000000000000000000000000000;
mem[658] = 64'b0101000111100000000000000000010000000000000000000000000000000000;
mem[659] = 64'b0101001010001000010001000000000001000001000000000000000000000000;
mem[660] = 64'b0101000111100000111001000101001010000000000010011100000000000000;
mem[661] = 64'b0101000111100000000000000000010000000000000000000000000000000000;
mem[662] = 64'b0101001011101000010001000000000001000001000000000000000000000000;
mem[663] = 64'b0101001100000000001000000000000000000001000000001000000000000010;
mem[664] = 64'b1001001100100000001000000000000000001000000000000000110000000000;
mem[665] = 64'b0101001101000000000000000000000000000001100000000100000000000010;
mem[666] = 64'b0101001101100000000000000000000000000100000000000000110000000010;
mem[667] = 64'b0101001110011000000000000000000000000001000000000100000000000010;
mem[668] = 64'b0101010010000000000000000000000010000000000000000000000000000000;
mem[669] = 64'b0101001111000000000000000000000000000001000000000000000000000000;
mem[670] = 64'b0101001111100000000000000000000000000001000000000000000000000000;
mem[671] = 64'b0101010000000000000000000000000000000001000000000000000000000000;
mem[672] = 64'b0101010000100000000000000000000000000001000000000000000000000000;
mem[673] = 64'b0101010001000000000000000000000000000001000000000000000000000000;
mem[674] = 64'b0101010001100000000000000000000000000001000000000000000000000000;
mem[675] = 64'b0101010010000000000000000000000000000001000000000000000000000000;
mem[676] = 64'b0101010010100000001001000000000000000001000000001000000000000010;
mem[677] = 64'b1001001100100000001001000000000000001000000000000000110000000000;
mem[678] = 64'b0101010011100000000000000000000000000100000000000000110000000010;
mem[679] = 64'b0101010100011000000000000000000000000001000000001100000000000010;
mem[680] = 64'b1001001100100000000000000000000000001000000000000000110000000000;
mem[681] = 64'b0101010101000000000000100000000000000001000000000100000100000000;
mem[682] = 64'b0101010101100000000000000000000000000100000000000000110000000000;
mem[683] = 64'b0101010110011000000000100000000000000001000000000100000100000000;
mem[684] = 64'b0101011010000000000000000000000010000000000000000000001000000000;
mem[685] = 64'b0101011010000000000000000000000010000000000000000000011000000000;
mem[686] = 64'b0101011010000000000000000000000010000000000000000000101000000000;
mem[687] = 64'b0101011010000000000000000000000010000000000000000000111000000000;
mem[688] = 64'b0101011010000000000000000000000010000000000000000000001000000000;
mem[689] = 64'b0101011010000000000000000000000010000000000000000000011000000000;
mem[690] = 64'b0101011010000000000000000000000010000000000000000000101000000000;
mem[691] = 64'b0101011010000000000000000000000010000000000000000000111000000000;
mem[692] = 64'b0101011010100000001010000000000000000001000000001000000000000000;
mem[693] = 64'b1001001100000000001010000000000000001000000000000000110000000000;
mem[694] = 64'b0101011100100000000000000000001000000000011010000000000000000000;
mem[695] = 64'b0101011111100000000000000000010000000000000100000000000000000000;
mem[696] = 64'b0101011100100000111001000101000000000000011000011100000000000000;
mem[697] = 64'b0101011101000000000000000000000000110000011000000000110000000000;
mem[698] = 64'b0101011101100000000000000000000000000100000000000000110000000001;
mem[699] = 64'b0101011110010010111001000101000000000000011101101100000000000000;
mem[700] = 64'b0101011110100000000000000000000000110000011100000000001000000000;
mem[701] = 64'b0101100000000000000000000000001000000010000000000000001000000001;
mem[702] = 64'b0101011011110010111001010101000000000000000011111100000000000000;
mem[703] = 64'b0101100000000000000000000000000000000001000000000000000000000000;
mem[704] = 64'b0101100000110010111001000101000000000001000001111100000000000000;
mem[705] = 64'b0101100010000000000000000000001000000000011010000000000000000000;
mem[706] = 64'b0101100101000000000000000000010000000000000100000000000000000000;
mem[707] = 64'b0101100010000000111001000101000000000000011000011100000000000000;
mem[708] = 64'b0101100010100000000000000000000000110000011000000000000000000000;
mem[709] = 64'b0101100011000010111001000011000000000000000001101100110000000000;
mem[710] = 64'b0101100011100000000000000000000000110100011100000000110000000000;
mem[711] = 64'b0101100100000010111001000011000000000000000001111100001000000000;
mem[712] = 64'b0101100101000000000000000000001000000010000000000000001000000000;
mem[713] = 64'b0101100001000000000000010000000000000000000010000000000000000000;
mem[714] = 64'b0101100101100000000000000000000000000001000000000000000000000000;
mem[715] = 64'b0101100110100000000000000000000000001000000000000000000000000001;
mem[716] = 64'b0101100110100000000000000000000000000100000000000000110000000001;
mem[717] = 64'b0101100111000000000000000000000000000000000000000000000010000001;
mem[718] = 64'b0101100111111011100011000000000000000000000000000000000010101101;
mem[719] = 64'b0101101000000000001011000000000000000001000000001100000000000000;
mem[720] = 64'b0101101001000000000000000000000000001000000000000000000000000000;
mem[721] = 64'b0101101001000000000000000000000000000100000000000000110000000000;
mem[722] = 64'b0101101001100000000000000000000000000000000000000000000010000000;
mem[723] = 64'b0101101010011011100011000000000000000000000000001100000011101100;
mem[724] = 64'b0101101010100000001011000000000000000001000000101100000000000000;
mem[725] = 64'b0101101011100000000000000000000000001000000000000000000000000001;
mem[726] = 64'b0101101011100000000000000000000000000100000000000000110000000001;
mem[727] = 64'b0101101100000000000000000000000000000000000000000000000010000001;
mem[728] = 64'b0101101100111011101011000000000000000000000000000000000010101101;
mem[729] = 64'b0101101101000000001011000000000000000001000000001100000000000000;
mem[730] = 64'b0101101110000000000000000000000000001000000000000000000000000000;
mem[731] = 64'b0101101110000000000000000000000000000100000000000000110000000000;
mem[732] = 64'b0101101110100000000000000000000000000000000000000000000010000000;
mem[733] = 64'b0101101111011011101011000000000000000000000000001100000011101100;
mem[734] = 64'b0101101111100000001011000000000000000001000000101100000000000000;
mem[735] = 64'b0101110000000011101001000000000000000001000000000100000000101100;
mem[736] = 64'b0101110000100000000000000000000000000100000000000000110000000000;
mem[737] = 64'b0101110001011011101001000000000000000001000000000100000000101100;
mem[738] = 64'b0101110001100001000001000001000000000001000000001000000000001110;
mem[739] = 64'b0101110010000000000000000000000000000100100000000000110000000010;
mem[740] = 64'b1001001100111001000001000001000000001000000000000000110000001110;
mem[741] = 64'b0101110011000010110001000001000000000001000000001000000000001110;
mem[742] = 64'b0101110011100000000000000000000000000100100000000000110000000010;
mem[743] = 64'b1001001100111010110001000001000000001000000000000000110000001110;
mem[744] = 64'b0101110100100000110000000000000000000001000000001000000000010010;
mem[745] = 64'b0101110101000000000000000000000000000100000000000000110000000010;
mem[746] = 64'b1001001100111000110000000000000000001000000000000000110000010010;
mem[747] = 64'b0101110110000000110000000000000000000001000000000100000000010010;
mem[748] = 64'b0101110110100000000000000000000000000100000000000000110000000010;
mem[749] = 64'b0101110111011000110000000000000000000001000000000100000000010010;
mem[750] = 64'b0101110111100000110001000000000000000001000000001100000000010010;
mem[751] = 64'b0101111000000000110001000000000000000001000000001000000000010010;
mem[752] = 64'b0101111000100000000000000000000000000100000000000000110000000010;
mem[753] = 64'b1001001100111000110001000000000000001000000000000000110000010010;
mem[754] = 64'b0101111010000000000000000000000000000000100000000000000000000000;
mem[755] = 64'b0101111010100000000000000000000000000000100000000000110000000000;
mem[756] = 64'b0101111010100000110001000000000000000001000000001000000000010000;
mem[757] = 64'b0101111011000000000000000000000000000100000000000000110000000000;
mem[758] = 64'b1001001100011000110001000000000000001000000000000000110000010000;
mem[759] = 64'b0101111100100000000000000000000000110000000000000000101000000000;
mem[760] = 64'b0101111110000000000000000000000000110000000000000000101000000000;
mem[761] = 64'b0101111101000000000000000000000000000100010000000000101000000000;
mem[762] = 64'b0101111101100000010001000011000000000000000001001100000000000000;
mem[763] = 64'b0101111110011000000000000000000000000001000000001000000000000000;
mem[764] = 64'b0101111110100000000000000000000000000100010000000000101000000000;
mem[765] = 64'b0101111111000000010001000011000000000000000001001100000000000000;
mem[766] = 64'b1001001100000000000000000000000000010000000000000000110000000000;
mem[767] = 64'b0110000000000000000000000000000000110000000000000000101000000000;
mem[768] = 64'b0110000000110000010001000011000000000100000001001100101000000000;
mem[769] = 64'b0110000001011000000000100000000000000001000000000000001100000000;
mem[770] = 64'b0110000001100000000000000000000000110000000000000000101000000000;
mem[771] = 64'b0110000010010000010001000011000000000100000001001100101000000000;
mem[772] = 64'b0110000010111000000000100000000000000001000000000000101100000000;
mem[773] = 64'b0110000011000000000000000000000000110000000000000000101000000000;
mem[774] = 64'b0110000011110000010001000011000000000100000001001100101000000000;
mem[775] = 64'b0110000100011000000000100000000000000001000000000000111100000000;
mem[776] = 64'b0110000100100000000000000000000000110000000000000000101000000000;
mem[777] = 64'b0110000101010000010001000011000000000100000001001100101000000000;
mem[778] = 64'b0110000101111000000000000000000000000001000000001100000000000000;
mem[779] = 64'b0110000110000000000000000000000000110000000000000000101000000000;
mem[780] = 64'b0110000110110000010001000011000000000100000001001100101000000000;
mem[781] = 64'b0110000111011000000000000000000000000001000000011100000000000000;
mem[782] = 64'b0110000111100000000000000000000000110000000000000000101000000000;
mem[783] = 64'b0110001000010000010001000011000000000100000001001100101000000000;
mem[784] = 64'b0110001000111000000000000000000000000001000000101100000000000000;
mem[785] = 64'b0110001001000000000000000000000000110000000000000000101000000000;
mem[786] = 64'b0110001001110000010001000011000000000100000001001100101000000000;
mem[787] = 64'b0110001010011000000000000000000000000001000000111100000000000000;
mem[788] = 64'b0110001010100000000000000000000000110000000000000000101000000000;
mem[789] = 64'b0110001011010000010001000011000000000100000001001100101000000000;
mem[790] = 64'b0110001011111000000000000000000000000001000001001100000000000000;
mem[791] = 64'b0110001100000000000000000000000000110000000000000000101000000000;
mem[792] = 64'b0110001100110000010001000011000000000100000001001100101000000000;
mem[793] = 64'b0110001101011000000000000000000000000001000001011100000000000000;
mem[794] = 64'b0110001101100000000000000000000000110000000000000000101000000000;
mem[795] = 64'b0110001110010000010001000011000000000100000001001100101000000000;
mem[796] = 64'b0110001110111000000000000000000000000001000001101100000000000000;
mem[797] = 64'b0110001111000000000000000000000000110000000000000000101000000000;
mem[798] = 64'b0110001111110000010001000011000000000100000001001100101000000000;
mem[799] = 64'b0110010000011000000000000000000000000001000001111100000000000000;
mem[800] = 64'b0110010000100000000000000000000000110000000000000000101000000000;
mem[801] = 64'b0110010001010000010001000011000000000100000001001100101000000000;
mem[802] = 64'b0110010001111001101000100000000000000001000000000000000000110000;
mem[803] = 64'b0110010010100000111001000011000000110000100001001100110000000000;
mem[804] = 64'b0110010011100000000000000000000000000100010000000000110000000000;
mem[805] = 64'b0110010011000000000000000000000000001000000000000000101000000000;
mem[806] = 64'b0110010011110000000000000000000000000011000000000000101000000000;
mem[807] = 64'b0110010100000000111001000011000000110000000001001100101000000000;
mem[808] = 64'b0110010100110000000000000000000000000011000000000000101000000000;
mem[809] = 64'b0110010101000000000000000000000000001000010000000000000000000000;
mem[810] = 64'b0110010101100000111001000011000000110000000001000000101000000000;
mem[811] = 64'b0110010110010000000000000000000000000011000001001100101000000000;
mem[812] = 64'b0110010110100000111001000011000000111000000001000000101000000000;
mem[813] = 64'b0110010111010000000000000000000000000011000001001100101000000000;
mem[814] = 64'b0110010111100000001010000000000000001000010000000000000000000000;
mem[815] = 64'b0110011000000000111001000011000000110000000001000000101000000000;
mem[816] = 64'b0110011000110000000000000000000000000011000001001100101000000000;
mem[817] = 64'b0110011001000000111001000011000000110000000001001100000000000000;
mem[818] = 64'b0110011001100000001001000000000000001000000000000000101000000000;
mem[819] = 64'b0110011010000000000000000000000000000011000000000000101000000000;
mem[820] = 64'b0110011010100000111001000011000000110000000001001100000000000000;
mem[821] = 64'b0110011011000000001001000000000000001000000000000000101000000000;
mem[822] = 64'b0110011011100000000000000000000000000011000000000000101000000000;
mem[823] = 64'b0110011100000000111001000011000000110000000001001100101000000000;
mem[824] = 64'b0110011100100000000000000000000000000011000000000000101000000000;
mem[825] = 64'b0110011101000000111001000011000000110000000000000000000000000000;
mem[826] = 64'b0110011101100000000000000000000000001000000000000000101000000000;
mem[827] = 64'b0110011110010000111001000011000000110010000100000000101000000000;
mem[828] = 64'b0110011110100000000000000000000000001000000000000000101000000000;
mem[829] = 64'b0110011111010000111001000011000000110010001000000000101000000000;
mem[830] = 64'b0110011111100000000000000000000000001000000000000000101000000000;
mem[831] = 64'b0110100000010000111001000011000000110010001100000000101000000000;
mem[832] = 64'b0110100000100000000000000000000000001000000000000000101000000000;
mem[833] = 64'b0110100001010000111001000011000000110010010000000000101000000000;
mem[834] = 64'b0110100001100000000000000000000000001000000000000000101000000000;
mem[835] = 64'b0110100010010000111001000011000000110010010100000000101000000000;
mem[836] = 64'b0110100010100000000000000000000000001000000000000000101000000000;
mem[837] = 64'b0110100011010000111001000011000000110010011000000000101000000000;
mem[838] = 64'b0110100011100000000000000000000000001000000000000000101000000000;
mem[839] = 64'b0110100100010000111001000011000000110010011100000000101000000000;
mem[840] = 64'b0110100100100000000000000000000000001000000000000000101000000000;
mem[841] = 64'b0110100101010000000000000000000000000011000001001100101000000000;
mem[842] = 64'b0110100101100000000000000000000000110000000000000000101000000000;
mem[843] = 64'b0110100110011000000000000000000000000100000001111100101000000000;
mem[844] = 64'b0110100110110000010001000011000000110000000000000000101000000000;
mem[845] = 64'b0110100111011000000000000000000000000100000001101100101000000000;
mem[846] = 64'b0110100111110000010001000011000000110000000000000000101000000000;
mem[847] = 64'b0110101000011000000000000000000000000100000001011100101000000000;
mem[848] = 64'b0110101000110000010001001001000000110000000000000000101000000000;
mem[849] = 64'b0110101001011000000000000000000000000100000000111100101000000000;
mem[850] = 64'b0110101001110000010001000011000000110000000000000000101000000000;
mem[851] = 64'b0110101010011000000000000000000000000100000000101100101000000000;
mem[852] = 64'b0110101010110000010001000011000000110000000000000000101000000000;
mem[853] = 64'b0110101011011000000000000000000000000100000000011100101000000000;
mem[854] = 64'b0110101011110000010001000011000000110000000000000000101000000000;
mem[855] = 64'b0110101100011000000000000000000000000100000000001100101000000000;
mem[856] = 64'b0110101100110000010001000011000000000001000001001100000000000000;
mem[857] = 64'b0110101101000010100001000101000000000001000000001000000000110110;
mem[858] = 64'b0110101101100000000000000000000000000100000000000000110000000010;
mem[859] = 64'b1001001100111010100001000101000000001000000000000000110000110110;
mem[860] = 64'b0110101110100000001000000000000010000000100000000000110010000010;
mem[861] = 64'b0110101111000010100000000000000000000001100000001000000011010110;
mem[862] = 64'b0110101111100000000000000000000000000100000010000000110000000010;
mem[863] = 64'b1001001100111010100000000000000000001000000000000000110011010110;
mem[864] = 64'b0110110000100010100001000000000000000001100000001000000011010110;
mem[865] = 64'b0110110001000000000000000000000000000100000000000000110000000010;
mem[866] = 64'b1001001100111010100001000000000000001000000000000000110011010110;
mem[867] = 64'b0110110000000000001001000000000010000000100000000000110010000000;
mem[868] = 64'b0110110010100010101001000101000000000001000000001000000000110110;
mem[869] = 64'b0110110011000000000000000000000000000100000000000000110000000010;
mem[870] = 64'b1001001100111010101001000101000000001000000000000000110000110110;
mem[871] = 64'b0110110100000000001000000000000010000000100000000000110010000010;
mem[872] = 64'b0110110100100010101000000000000000000001100000001000000011010110;
mem[873] = 64'b0110110101000000000000000000000000000100000010000000110000000010;
mem[874] = 64'b1001001100111010101000000000000000001000000000000000110011010110;
mem[875] = 64'b0110110110000010101001000000000000000001100000001000000011010110;
mem[876] = 64'b0110110110100000000000000000000000000100000000000000110000000010;
mem[877] = 64'b1001001100111010101001000000000000001000000000000000110011010110;
mem[878] = 64'b0110110101100000001001000000000010000000100000000000110010000000;
mem[879] = 64'b0110111000000000000000000000000000110000000000000000101000000000;
mem[880] = 64'b0110111000110000010001000011000000000100000001001100101000000000;
mem[881] = 64'b0110111001011000000000000000000001000001000000000000000000000000;
mem[882] = 64'b0110111001100000000000000000000000110000000000000000101000000000;
mem[883] = 64'b0110111010010000010001000011000000000100000001001100101000000000;
mem[884] = 64'b0110111010111000000000000000000001000000010000000000000000000000;
mem[885] = 64'b0110111011000000010001000000000000000001000001001100000000000000;
mem[886] = 64'b0110111011100000000000000000000000110000000000000000101000000000;
mem[887] = 64'b0110111100010000010001000011000000110100000000000000101000000000;
mem[888] = 64'b0110111100111000000000000000000001000000000000000000101000000000;
mem[889] = 64'b0110111101010000010001000011000000000100000001001100101000000000;
mem[890] = 64'b0110111101111000000000000000000000000001000000000000011100000000;
mem[891] = 64'b0110111110000000000000000000000000110000000000000000101000000000;
mem[892] = 64'b0110111110110000010001000011000000110100000000000000101000000000;
mem[893] = 64'b0110111111011000000000000000000001000000000000000000101000000000;
mem[894] = 64'b0110111111110000010001000011000000110100000000000000101000000000;
mem[895] = 64'b0111000000010000010001000000000000000000000001001100000000000000;
mem[896] = 64'b0111000000111000000000000000000000000001000000000000011100000000;
mem[897] = 64'b0111000001000000000000000000000000110000000000000000101000000000;
mem[898] = 64'b0111000001110000010001000011000000110100000000000000101000000000;
mem[899] = 64'b0111000010011000000000000000000001000000000000000000101000000000;
mem[900] = 64'b0111000010100000000000000000000000000100000000000000101000000000;
mem[901] = 64'b0111000011011000000000000000000000000000000000000000011100000000;
mem[902] = 64'b0111000011110000010001000011000000110000000000000000101000000000;
mem[903] = 64'b0111000100011001101000000000000000000100000000000000101000110000;
mem[904] = 64'b0111000100110000010001100011000000000001000001001100000000000000;
mem[905] = 64'b0111000101000010011001000101000000000001000000001000000000110110;
mem[906] = 64'b0111000101100000000000000000000000000100000000000000110000000010;
mem[907] = 64'b1001001100111010011001000101000000001000000000000000110000110110;
mem[908] = 64'b0111000110100000001000000000000010000000100000000000110010000010;
mem[909] = 64'b0111000111000010011000000000000000000001100000001000000011010110;
mem[910] = 64'b0111000111100000000000000000000000000100000010000000110000000010;
mem[911] = 64'b1001001100111010011000000000000000001000000000000000110011010110;
mem[912] = 64'b0111001000100010011001000000000000000001100000001000000011010110;
mem[913] = 64'b0111001001000000000000000000000000000100000000000000110000000010;
mem[914] = 64'b1001001100111010011001000000000000001000000000000000110011010110;
mem[915] = 64'b0111001000000000001001000000000010000000100000000000110010000000;
mem[916] = 64'b0111001010100010010001000101000000000001000000001000000000110110;
mem[917] = 64'b0111001011000000000000000000000000000100000000000000110000000010;
mem[918] = 64'b1001001100111010010001000101000000001000000000000000110000110110;
mem[919] = 64'b0111001100000000001000000000000010000000100000000000110010000010;
mem[920] = 64'b0111001100100010010000000000000000000001100000001000000011010110;
mem[921] = 64'b0111001101000000000000000000000000000100000010000000110000000010;
mem[922] = 64'b1001001100111010010000000000000000001000000000000000110011010110;
mem[923] = 64'b0111001110000010010001000000000000000001100000001000000011010110;
mem[924] = 64'b0111001110100000000000000000000000000100000000000000110000000010;
mem[925] = 64'b1001001100111010010001000000000000001000000000000000110011010110;
mem[926] = 64'b0111001101100000001001000000000010000000100000000000110010000000;
mem[927] = 64'b0111010000000010001001000101000000000001000000001000000000010010;
mem[928] = 64'b0111010000100000000000000000000000000100000000000000110000000010;
mem[929] = 64'b1001001100111010001001000101000000001000000000000000110000010010;
mem[930] = 64'b0111010001100000001000000000000010000000100000000000110010000010;
mem[931] = 64'b0111010010000010001000000000000000000001100000001000000011111010;
mem[932] = 64'b0111010010100000000000000000000000000100000010000000110000000010;
mem[933] = 64'b1001001100111010001000000000000000001000000000000000110011111010;
mem[934] = 64'b0111010011100010001001000000000000000001100000001000000011111010;
mem[935] = 64'b0111010100000000000000000000000000000100000000000000110000000010;
mem[936] = 64'b1001001100111010001001000000000000001000000000000000110011111010;
mem[937] = 64'b0111010011000000001001000000000010000000100000000000110010000000;
mem[938] = 64'b0111010101100001001000000000000000000001000000001000000000001110;
mem[939] = 64'b0111010110000000000000000000000000000100000000000000110000000010;
mem[940] = 64'b1001001100111001001000000000000000001000000000000000110000001110;
mem[941] = 64'b0111010111000001010000000000000000000001000000000100000000001110;
mem[942] = 64'b0111010111100000000000000000000000000100000000000000110000000010;
mem[943] = 64'b0111011000011001010000000000000000000001000000000100000000001110;
mem[944] = 64'b0111011000100001001001000000000000000001000000001100000000001110;
mem[945] = 64'b0111011001000001001001000000000000000001000000001000000000001110;
mem[946] = 64'b0111011001100000000000000000000000000100000000000000110000000010;
mem[947] = 64'b1001001100111001001001000000000000001000000000000000110000001110;
mem[948] = 64'b0111011011000000000000000000000000000000100000000000000000000000;
mem[949] = 64'b0111011011100000000000000000000000000000100000000000110000000000;
mem[950] = 64'b0111011011100001001001000000000000000001000000001000000000001100;
mem[951] = 64'b0111011100000000000000000000000000000100000000000000110000000000;
mem[952] = 64'b1001001100011001001001000000000000001000000000000000110000001100;
mem[953] = 64'b0111011110000000000000000000001000110000011110000000000000000000;
mem[954] = 64'b0111011111100000000000000000010000000000000100000000000000000000;
mem[955] = 64'b0111011110000000111001000101000000000000011100011100001000000000;
mem[956] = 64'b0111011110100000000000000000000000000100000000000000001010000001;
mem[957] = 64'b0111100000011001000011000000001000000000000000000000000000001101;
mem[958] = 64'b0111011101010010111001010101001100110000000011111100001000000000;
mem[959] = 64'b0111100000000000000000000000000000000001000000000000000000000000;
mem[960] = 64'b0111100000110010111001000101000000000001000001111100000000000000;
mem[961] = 64'b0111100010000000000000000000001000110000011110000000000000000000;
mem[962] = 64'b0111100011100000000000000000010000000000000100000000000000000000;
mem[963] = 64'b0111100010000000111001000101000000000000011100011100001000000000;
mem[964] = 64'b0111100010100000000000000000000000000100000000000000001010000000;
mem[965] = 64'b0111100100011001000011000000001000000000000000000000000000001100;
mem[966] = 64'b0111100001010010111001010011001100110000000011111100001000000000;
mem[967] = 64'b0111100100000000000000000000000000000001000000000000000000000000;
mem[968] = 64'b0111100100110010111001000011000000000001000001111100000000000000;
mem[969] = 64'b0111100101000010000001000101000000000001000000001000000000010010;
mem[970] = 64'b0111100101100000000000000000000000000100000000000000110000000010;
mem[971] = 64'b1001001100111010000001000101000000001000000000000000110000010010;
mem[972] = 64'b0111100110100000001000000000000010000000100000000000110010000010;
mem[973] = 64'b0111100111000010000000000000000000000001100000001000000011111010;
mem[974] = 64'b0111100111100000000000000000000000000100000010000000110000000010;
mem[975] = 64'b1001001100111010000000000000000000001000000000000000110011111010;
mem[976] = 64'b0111101000100010000001000000000000000001100000001000000011111010;
mem[977] = 64'b0111101001000000000000000000000000000100000000000000110000000010;
mem[978] = 64'b1001001100111010000001000000000000001000000000000000110011111010;
mem[979] = 64'b0111101000000000001001000000000010000000100000000000110010000000;
mem[980] = 64'b0111101010100001111001000101000000000001000000001000000000010010;
mem[981] = 64'b0111101011000000000000000000000000000100000000000000110000000010;
mem[982] = 64'b1001001100111001111001000101000000001000000000000000110000010010;
mem[983] = 64'b0111101100000000001000000000000010000000100000000000110010000010;
mem[984] = 64'b0111101100100001111000000000000000000001100000001000000011111010;
mem[985] = 64'b0111101101000000000000000000000000000100000010000000110000000010;
mem[986] = 64'b1001001100111001111000000000000000001000000000000000110011111010;
mem[987] = 64'b0111101110000001111001000000000000000001100000001000000011111010;
mem[988] = 64'b0111101110100000000000000000000000000100000000000000110000000010;
mem[989] = 64'b1001001100111001111001000000000000001000000000000000110011111010;
mem[990] = 64'b0111101101100000001001000000000010000000100000000000110010000000;
mem[991] = 64'b0111110000000000000000000000000000001000000000000000000000000001;
mem[992] = 64'b0111110001100000000000000000001000000000011110000000000000000000;
mem[993] = 64'b0111110100100000000000000000010000000000000100000000000000000000;
mem[994] = 64'b0111110001100000111001000101000000000000011100011100000000000000;
mem[995] = 64'b0111110010000000000000000000000000110000011100000000000000000000;
mem[996] = 64'b0111110010100010111001000101000000000000000001111100000000000000;
mem[997] = 64'b0111110011000000000000000000000000000000000000000000000000000001;
mem[998] = 64'b0111110011100000000000000000000000001000000000000000001000000001;
mem[999] = 64'b0111110100100000000000000000001000000010000000000000001000000001;
mem[1000] = 64'b0111110000100000000000010000000000000000000010000000000000000000;
mem[1001] = 64'b0111110101000000000000000000000000000001000000000000000000000000;
mem[1002] = 64'b0111110110100000000000000000001000001000011110000000000000000000;
mem[1003] = 64'b0111111000100000000000000000010000000000000100000000000000000000;
mem[1004] = 64'b0111110110100000111001000101000000000000011100011100000000000000;
mem[1005] = 64'b0111110111000000000000000000000000110000011100000000000000000000;
mem[1006] = 64'b0111110111100010111001000011000000000000000001111100001000000000;
mem[1007] = 64'b0111111000100000000000000000001000000010000000000000001000000000;
mem[1008] = 64'b0111110101100000000000010000000000000000000010000000000000000000;
mem[1009] = 64'b0111111001000000000000000000000000000001000000000000000000000000;
mem[1010] = 64'b0111111001100000111000000000000000000001000000001000000000001110;
mem[1011] = 64'b0111111010000000000000000000000000000100000000000000110000000010;
mem[1012] = 64'b1001001100111000111000000000000000001000000000000000110000001110;
mem[1013] = 64'b0111111011000001000000000000000000000001000000000100000000001110;
mem[1014] = 64'b0111111011100000000000000000000000000100000000000000110000000010;
mem[1015] = 64'b0111111100011001000000000000000000000001000000000100000000001110;
mem[1016] = 64'b0111111100100000111001000000000000000001000000001100000000001110;
mem[1017] = 64'b0111111101000000111001000000000000000001000000001000000000001110;
mem[1018] = 64'b0111111101100000000000000000000000000100000000000000110000000010;
mem[1019] = 64'b1001001100111000111001000000000000001000000000000000110000001110;
mem[1020] = 64'b0111111111000000000000000000000000000000100000000000000000000000;
mem[1021] = 64'b0111111111100000000000000000000000000000100000000000110000000000;
mem[1022] = 64'b0111111111100000111001000000000000000001000000001000000000001100;
mem[1023] = 64'b1000000000000000000000000000000000000100000000000000110000000000;
mem[1024] = 64'b1001001100011000111001000000000000001000000000000000110000001100;
mem[1025] = 64'b1000000001000000100000000000000000000001000000000000000000010010;
mem[1026] = 64'b1000000001100000000000000000000000000100000000000000110000000010;
mem[1027] = 64'b1000000010011000100000000000000000000001000000000000000000010010;
mem[1028] = 64'b1000000010100000100001000000000000000001000000000000000000010010;
mem[1029] = 64'b1000000011000000100001000000000000000001000000000000000000010001;
mem[1030] = 64'b1000000011100000000000000000000000000100000000000000110000000001;
mem[1031] = 64'b1000000100011000100001000000000000000001000000000000000000010001;
mem[1032] = 64'b1000000100100000100001000000000000000001000000000000000000010000;
mem[1033] = 64'b1000000101000000000000000000000000000100000000000000110000000000;
mem[1034] = 64'b1000000101111000100001000000000000000001000000000000000000010000;
mem[1035] = 64'b1000001000000000000000000000000000110000000000000000000000000010;
mem[1036] = 64'b1000000110100000000000000000000000000100000000000000110000000010;
mem[1037] = 64'b1000000111000000001000000000000000110000000000000000000000000010;
mem[1038] = 64'b1000000111111000000000000000000000000000000000000100000000000010;
mem[1039] = 64'b1001001100110000000000000000000000011000000000000000110000000010;
mem[1040] = 64'b1000001000100000001000000000000000000000000000001000000000000010;
mem[1041] = 64'b1000001001010000000000000000000000000001000000000100000000000010;
mem[1042] = 64'b1000001001100000000000000000000000110000000000000000000000000000;
mem[1043] = 64'b1000001010000000000000000000000000000000000000011100000000000000;
mem[1044] = 64'b1000001010110000000000000000000000000001000000001100000000000000;
mem[1045] = 64'b1000001011000000000000000000000000110000000000000000000000000000;
mem[1046] = 64'b1000001011100000000000000000000000000000000000101100000000000000;
mem[1047] = 64'b1000001100010000000000000000000000000001000000001100000000000000;
mem[1048] = 64'b1000001100100000000000000000000000110000000000000000000000000000;
mem[1049] = 64'b1000001101000000000000000000000000000000000000111100000000000000;
mem[1050] = 64'b1000001101110000000000000000000000000001000000001100000000000000;
mem[1051] = 64'b1000001110000000000000000000000000110000000000000000000000000000;
mem[1052] = 64'b1000001110100000000000000000000000000000000001001100000000000000;
mem[1053] = 64'b1000001111010000000000000000000000000001000000001100000000000000;
mem[1054] = 64'b1000001111100000000000000000000000110000000000000000000000000000;
mem[1055] = 64'b1000010000000000000000000000000000000000000001011100000000000000;
mem[1056] = 64'b1000010000110000000000000000000000000001000000001100000000000000;
mem[1057] = 64'b1000010001000000000000000000000000110000000000000000000000000000;
mem[1058] = 64'b1000010001100000000000000000000000000000000001101100000000000000;
mem[1059] = 64'b1000010010010000000000000000000000000001000000001100000000000000;
mem[1060] = 64'b1000010010100000000000000000000000110000000000000000000000000000;
mem[1061] = 64'b1000010011000000000000000000000000000000000001111100000000000000;
mem[1062] = 64'b1000010011110000000000000000000000000001000000001100000000000000;
mem[1063] = 64'b1000010100000000000000000000000000000000001100000000000010000000;
mem[1064] = 64'b1000010100100000000000000000000000110000000000000000000000000000;
mem[1065] = 64'b1000010101010000010011000000000000110000000000000000110000000000;
mem[1066] = 64'b1000010101111000000000000000000000000101000000001100110000000001;
mem[1067] = 64'b1000010110000000101000000000000000000001000000001000000000010010;
mem[1068] = 64'b1000010110100000000000000000000000000100000000000000110000000010;
mem[1069] = 64'b1001001100111000101000000000000000001000000000000000110000010010;
mem[1070] = 64'b1000010111100000101000000000000000000001000000000100000000010010;
mem[1071] = 64'b1000011000000000000000000000000000000100000000000000110000000010;
mem[1072] = 64'b1000011000111000101000000000000000000001000000000100000000010010;
mem[1073] = 64'b1000011001000000101001000000000000000001000000001100000000010010;
mem[1074] = 64'b1000011001100000101001000000000000000001000000001000000000010010;
mem[1075] = 64'b1000011010000000000000000000000000000100000000000000110000000010;
mem[1076] = 64'b1001001100111000101001000000000000001000000000000000110000010010;
mem[1077] = 64'b1000011011100000000000000000000000000000100000000000000000000000;
mem[1078] = 64'b1000011100000000000000000000000000000000100000000000110000000000;
mem[1079] = 64'b1000011100000000101001000000000000000001000000001000000000010000;
mem[1080] = 64'b1000011100100000000000000000000000000100000000000000110000000000;
mem[1081] = 64'b1001001100011000101001000000000000001000000000000000110000010000;
mem[1082] = 64'b0010010110100000001001000010000000000000000000000000000010000000;
mem[1083] = 64'b0010100110000000000000000000000010000000100000000000110000000010;
mem[1084] = 64'b0101110111100000000000000000000010000000100000000000110000000010;
mem[1085] = 64'b0010011110100000000000000000000010000000100000000000110000000010;
mem[1086] = 64'b0111011000100000000000000000000010000000100000000000110000000010;
mem[1087] = 64'b0010101101100000000000000000000010000000100000000000110000000010;
mem[1088] = 64'b0111111100100000000000000000000010000000100000000000110000000010;
mem[1089] = 64'b1000011001000000000000000000000010000000100000000000110000000010;
mem[1090] = 64'b0011001001100000000000000000000010000000100000000000110000000010;
mem[1091] = 64'b0010100111100000000000000000000010000000000000000000110000000000;
mem[1092] = 64'b0101111001000000000000000000000010000000000000000000110000000000;
mem[1093] = 64'b0010100000000000000000000000000010000000000000000000110000000000;
mem[1094] = 64'b0111011010000000000000000000000010000000000000000000110000000000;
mem[1095] = 64'b0010101111000000000000000000000010000000000000000000110000000000;
mem[1096] = 64'b0111111110000000000000000000000010000000000000000000110000000000;
mem[1097] = 64'b1000011010100000000000000000000010000000000000000000110000000000;
mem[1098] = 64'b0011001011000000000000000000000010000000000000000000110000000000;
mem[1099] = 64'b0101111011100000000000000000000010000000010000000000000000000000;
mem[1100] = 64'b1000100110100000000000000000000000000001000000000000000000000000;
mem[1101] = 64'b1000100111000000000000000000000000000001000000000000000000000000;
mem[1102] = 64'b1000100111100000000000000000000000000001000000000000000000000000;
mem[1103] = 64'b1000101000000000000000000000000000000001000000000000000000000000;
mem[1104] = 64'b1000101000100000000000000000000000000001000000000000000000000000;
mem[1105] = 64'b1000101001000000000000000000000000000001000000000000000000000000;
mem[1106] = 64'b1000101001100000000000000000000000000001000000000000000000000000;
mem[1107] = 64'b0111000100100000000000000000000010000000100000000000110000000010;
mem[1108] = 64'b0111001010000000000000000000000010000000100000000000110000000010;
mem[1109] = 64'b0110101100100000000000000000000010000000100000000000110000000010;
mem[1110] = 64'b0110110010000000000000000000000010000000100000000000110000000010;
mem[1111] = 64'b0111100100100000000000000000000010000000100000000000110000000010;
mem[1112] = 64'b0111101010000000000000000000000010000000100000000000110000000010;
mem[1113] = 64'b0111100100100000000000000000000010000000100000000000110000000010;
mem[1114] = 64'b0111001111100000000000000000000010000000100000000000110000000010;
mem[1115] = 64'b0111001000000000001001000000000010000000100000000000110010000001;
mem[1116] = 64'b0111001101100000001001000000000010000000100000000000110010000001;
mem[1117] = 64'b0110110000000000001001000000000010000000100000000000110010000001;
mem[1118] = 64'b0110110101100000001001000000000010000000100000000000110010000001;
mem[1119] = 64'b0111101000000000001001000000000010000000100000000000110010000001;
mem[1120] = 64'b0111101101100000001001000000000010000000100000000000110010000001;
mem[1121] = 64'b0111101000000000001001000000000010000000100000000000110010000001;
mem[1122] = 64'b0111010011000000001001000000000010000000100000000000110010000001;
mem[1123] = 64'b0111001001100000001001000000000000000000000000000000000010000001;
mem[1124] = 64'b0111001111000000001001000000000000000000000000000000000010000001;
mem[1125] = 64'b0110110001100000001001000000000000000000000000000000000010000001;
mem[1126] = 64'b0110110111000000001001000000000000000000000000000000000010000001;
mem[1127] = 64'b0111101001100000001001000000000000000000000000000000000010000001;
mem[1128] = 64'b0111101111000000001001000000000000000000000000000000000010000001;
mem[1129] = 64'b0111101001100000001001000000000000000000000000000000000010000001;
mem[1130] = 64'b0111010100100000001001000000000000000000000000000000000010000001;
mem[1131] = 64'b0111000110000000000000000000000000000000100010000000110000000010;
mem[1132] = 64'b0111001011100000000000000000000000000000100010000000110000000010;
mem[1133] = 64'b0110101110000000000000000000000000000000100010000000110000000010;
mem[1134] = 64'b0110110011100000000000000000000000000000100010000000110000000010;
mem[1135] = 64'b0111100110000000000000000000000000000000100010000000110000000010;
mem[1136] = 64'b0111101011100000000000000000000000000000100010000000110000000010;
mem[1137] = 64'b0111100110000000000000000000000000000000100010000000110000000010;
mem[1138] = 64'b0111010001000000000000000000000000000000100010000000110000000010;
mem[1139] = 64'b1000000010100000000000000000000010000000100000000000110000000001;
mem[1140] = 64'b1000000010100000000000000000000010000000100000000000110000000001;
mem[1141] = 64'b0101110010100000000000000000000010000000100000000000110000000001;
mem[1142] = 64'b0101110001000000000000000000000010000000100000000000110000000001;
mem[1143] = 64'b0101100101100000000000000000000010000000100000000000110000000001;
mem[1144] = 64'b0101101010100000000000000000000010000000100000000000110000000001;
mem[1145] = 64'b0011011001000000000000000000000010000000100000000000110000000001;
mem[1146] = 64'b0011011111100000000000000000000010000000100000000000110000000001;
mem[1147] = 64'b1000000100000000000000000000000010000000100000000000110000000000;
mem[1148] = 64'b1000000100000000000000000000000010000000100000000000110000000000;
mem[1149] = 64'b0101110010100000000000000000000010000000100000000000110000000000;
mem[1150] = 64'b0101110001000000000000000000000010000000100000000000110000000000;
mem[1151] = 64'b0101101000000000000000000000000010000000100000000000110000000000;
mem[1152] = 64'b0101101101000000000000000000000010000000100000000000110000000000;
mem[1153] = 64'b0011011100100000000000000000000010000000100000000000110000000000;
mem[1154] = 64'b0011100010000000000000000000000010000000100000000000110000000000;
mem[1155] = 64'b0011111000000000000000000000000010000000100000000000110000000000;
mem[1156] = 64'b0011111001100000000000000000000010000000100000000000110000000000;
mem[1157] = 64'b0010111001000000000000000000000010000000100000000000110000000000;
mem[1158] = 64'b0010111111100000000000000000000010000000000000000000011000000000;
mem[1159] = 64'b0100101101100000000000000000000010000000100000000000110000000000;
mem[1160] = 64'b0100101111000000000000000000000010000000100000000000110000000000;
mem[1161] = 64'b0110010001100000000000000000000010000000010000000000110000000000;
mem[1162] = 64'b1000011101000000000000000000000000000000000000000000000000000000;
mem[1163] = 64'b1001000110000000001001000001000000000000000000001100000000000000;
mem[1164] = 64'b1001000110100000001001000001000000000000000000011100000000000000;
mem[1165] = 64'b1001000111000000001001000001000000000000000000101100000000000000;
mem[1166] = 64'b1001000111100000001001000001000000000000000000111100000000000000;
mem[1167] = 64'b1001001000000000001001000001000000000000000001001100000000000000;
mem[1168] = 64'b1001001000100000001001000001000000000000000001011100000000000000;
mem[1169] = 64'b1001001001000000001001000001000000000000000001101100000000000000;
mem[1170] = 64'b1001001001100000001001000001000000000000000001111100000000000000;
mem[1171] = 64'b1001001010000000001001000001000000000000000000000000001100000000;
mem[1172] = 64'b1001001010100000001001000110000000000000000000000000011100000000;
mem[1173] = 64'b1001001011000000001001000001000000000000000000000000101100000000;
mem[1174] = 64'b1001001011100000001001000001000000000000000000000000111100000000;
mem[1175] = 64'b0010000000000000000000000000000000000001000000000000000000000000;
mem[1176] = 64'b1001001100100000000000000000000000000011000000000000110000000000;
mem[1177] = 64'b1001001101000000000000000000000000000011000000000000110000000010;
mem[1178] = 64'b0010000001000000000000000000000000000000000000000000000010000000;
mem[1179] = 64'b0010000001000000001010000000000000000000000000000000000010000000;
mem[1180] = 64'b1001001110100000000000000000000000000100000000000000111000000001;
mem[1181] = 64'b1001001111011000000000000000000000000000000000000000000010000000;
mem[1182] = 64'b0010000001010000010001000101000000110000000000000000000000000000;
mem[1183] = 64'b1001010000000000000000000000000000000100000000000000111000000000;
mem[1184] = 64'b1001010000111000000000000000000000000000000000000000000010000000;
mem[1185] = 64'b0010000001010000010001000011000000110000000000000000000000000000;
mem[1186] = 64'b1001010001100000000000000000000000000010000000000000111000000001;
mem[1187] = 64'b0010000001010000010001000101000000110000000000000000000000000000;
mem[1188] = 64'b1001010010100000000000000000000000000010000000000000111000000000;
mem[1189] = 64'b0010000001010000010001000011000000110000000000000000000000000000;
mem[1190] = 64'b1001010011100000000000000000100000000100000000000000111000000001;
mem[1191] = 64'b0010000001011000000000000000000000000000000000000000000010000000;
mem[1192] = 64'b1001010100100000000000000000100000000100000000000000111000000000;
mem[1193] = 64'b0010000001011000000000000000000000000000000000000000000010000000;
mem[1194] = 64'b0010000001000000000000000000100000000010000000000000111000000001;
mem[1195] = 64'b0010000001000000000000000000100000000010000000000000111000000000;	
end

always_comb begin
    case (current.immediate)
    1: microcode_immediate = 16'h0;
    2: microcode_immediate = 16'h18;
    3: microcode_immediate = 16'h2;
    4: microcode_immediate = 16'h14;
    5: microcode_immediate = 16'h1;
    6: microcode_immediate = 16'hffff;
    7: microcode_immediate = 16'hc;
    8: microcode_immediate = 16'hff;
    9: microcode_immediate = 16'h4;
    10: microcode_immediate = 16'h10;
    11: microcode_immediate = 16'h8;
    default: microcode_immediate = 16'h0;
    endcase
end

always_comb begin
    case (current.update_flags)
    0: update_flags = 9'h0;
    1: update_flags = 9'h5;
    2: update_flags = 9'h1a;
    3: update_flags = 9'h11f;
    4: update_flags = 9'h11b;
    5: update_flags = 9'h1;
    6: update_flags = 9'h1f;
    7: update_flags = 9'h40;
    8: update_flags = 9'h80;
    9: update_flags = 9'h11e;
    10: update_flags = 9'h60;
    11: update_flags = 9'h109;
    12: update_flags = 9'h1ff;
    13: update_flags = 9'h101;
    14: update_flags = 9'h1b;
    default: update_flags = 9'h0;
    endcase
end

assign a_sel = current.a_sel;
assign alu_op = current.alu_op;
assign b_sel = current.b_sel;
assign ext_int_yield = current.ext_int_yield;
assign io = current.io;
assign load_ip = current.load_ip;
assign mar_wr_sel = current.mar_wr_sel;
assign mar_write = current.mar_write;
assign mdr_write = current.mdr_write;
assign mem_read = current.mem_read;
assign mem_write = current.mem_write;
assign next_instruction = current.next_instruction;
assign ra_modrm_rm_reg = current.ra_modrm_rm_reg;
assign ra_sel = current.ra_sel;
assign rb_cl = current.rb_cl;
assign rd_sel = current.rd_sel;
assign rd_sel_source = current.rd_sel_source;
assign reg_wr_source = current.reg_wr_source;
assign segment = current.segment;
assign segment_force = current.segment_force;
assign segment_wr_en = current.segment_wr_en;
assign tmp_wr_en = current.tmp_wr_en;
assign tmp_wr_sel = current.tmp_wr_sel;

assign fifo_rd_en = starting_instruction;
assign starting_instruction = !stall && (next_addr == {{addr_bits-8{1'b0}}, next_instruction_value.opcode});
assign modrm_start = addr == modrm_wait_address ||
    (addr == next_instruction_address && !fifo_empty && next_instruction_value.has_modrm);
wire has_rep_prefix = cur_instruction.rep != REP_PREFIX_NONE;
reg rep_complete;
assign debug_stopped = addr == debug_wait_address;
assign multibit_shift = cur_instruction.opcode == 8'hd2 ||
                        cur_instruction.opcode == 8'hd3 ||
                        cur_instruction.opcode == 8'hc0 ||
                        cur_instruction.opcode == 8'hc1;
assign do_escape_fault = cur_instruction.opcode[7:3] == 5'b11011 && next_addr == do_int_address;
reg nmi_pending;
reg ext_int_inhibit;
wire take_nmi = (nmi_pending | nmi_pulse) & !ext_int_inhibit & !current.ext_int_inhibit;
wire take_irq = intr & int_enabled & !ext_int_inhibit & !current.ext_int_inhibit;
wire do_single_step = current.next_instruction & !ext_int_inhibit &
    trap_flag_set & current.next != debug_wait_address & !current.ext_int_inhibit;
assign start_interrupt = next_addr == nmi_address ||
                         next_addr == irq_address;
assign irq_to_mdr = next_addr == irq_address;
reg trap_flag_set;
assign is_hlt = cur_instruction.opcode == 8'hf4;
reg seized;
wire seizing = debug_seize & ~seized;
assign loop_next = !stall && current.jump_type == JumpType_LOOP_DONE;
assign reg_wr_en = current.rd_sel_source != RDSelSource_NONE & ~segment_wr_en;
assign next_microinstruction = addr != next_addr;
assign lock = cur_instruction.lock;

always_comb begin
    case (current.width)
    WidthType_W8: width = 1'b1;
    WidthType_W16: width = 1'b0;
    WidthType_WAUTO: width = ~cur_instruction.opcode[0];
    default: width = 1'b0;
    endcase
end

always_ff @(posedge clk)
    inta <= next_addr == irq_address && addr != irq_address;

always_ff @(posedge clk or posedge reset)
    if (reset)
        trap_flag_set <= 1'b0;
    else if (next_addr == single_step_address)
        trap_flag_set <= 1'b0;
    else if (starting_instruction)
        trap_flag_set <= tf;

always_ff @(posedge clk or posedge reset)
    if (reset)
        ext_int_inhibit <= 1'b0;
    else if (current.ext_int_inhibit && current.next != debug_wait_address)
        ext_int_inhibit <= 1'b1;
    else if (starting_instruction && !stall)
        ext_int_inhibit <= 1'b0;

//`ifdef verilator
//initial $readmemh({"microcode.hex"}, mem);
//`endif

always_comb begin
    case (cur_instruction.rep)
    REP_PREFIX_E: rep_complete = ~zf;
    REP_PREFIX_NE: rep_complete = zf;
    default: rep_complete = 1'b0;
    endcase
end

always_ff @(posedge clk or posedge reset)
    if (reset)
        nmi_pending <= 1'b0;
    else if (next_addr == nmi_address)
        nmi_pending <= 1'b0;
    else if (nmi_pulse)
        nmi_pending <= 1'b1;

always_ff @(posedge clk or posedge reset)
    if (reset)
        seized <= 1'b0;
    else if (debug_stopped)
        seized <= 1'b1;
    else if (!debug_seize)
        seized <= 1'b0;

always_comb begin
    unique case (current.jump_type)
    JumpType_RM_REG_MEM: jump_target = current.next + {{addr_bits-1{1'b0}}, ~rm_is_reg};
    JumpType_OPCODE: jump_target = !fifo_empty ? {{addr_bits-8{1'b0}}, next_instruction_value.opcode} : addr;
    JumpType_DISPATCH_REG: jump_target = current.next + {{addr_bits-3{1'b0}}, modrm_reg};
    JumpType_HAS_NO_REP_PREFIX: jump_target = ~has_rep_prefix ? current.next : addr + 1'b1;
    JumpType_ZERO: jump_target = zf ? current.next : addr + 1'b1;
    JumpType_REP_NOT_COMPLETE: jump_target = !rep_complete ? current.next : addr + 1'b1;
    JumpType_RB_ZERO: jump_target = rb_zero ? current.next : addr + 1'b1;
    JumpType_LOOP_DONE: jump_target = loop_done ? current.next : addr + 1'b1;
    JumpType_JUMP_TAKEN: jump_target = jump_taken ? current.next : addr + 1'b1;
    default: jump_target = current.next;
    endcase
end

always_comb begin
    if (reset)
        next_addr = reset_address;
    else if (debug_stopped && debug_run)
        next_addr = {{addr_bits - 9{1'b0}}, 1'b1, debug_addr};
    else if (stall)
        next_addr = addr;
    else if (current.ext_int_yield && seizing)
        next_addr = debug_wait_address;
    else if (current.ext_int_yield && take_nmi)
        next_addr = nmi_address;
    else if (current.ext_int_yield && take_irq)
        next_addr = irq_address;
    else if (addr == next_instruction_address && !fifo_empty && !fifo_resetting &&
             next_instruction_value.invalid)
        next_addr = bad_opcode_address;
    else if (current.jump_type != JumpType_UNCONDITIONAL)
        next_addr = jump_target;
    else if (divide_error)
        next_addr = divide_error_address;
    else if (current.next_instruction && take_nmi)
        next_addr = nmi_address;
    else if (current.next_instruction && take_irq)
        next_addr = irq_address;
    else if ((current.next_instruction && do_single_step) ||
             (is_hlt && trap_flag_set))
        next_addr = single_step_address;
    else if (current.next_instruction && debug_seize)
        next_addr = debug_wait_address;
    else if (current.next_instruction || (is_hlt && intr))
        next_addr = !fifo_empty && !fifo_resetting ?
            (next_instruction_value.has_modrm ? modrm_wait_address :
             {{addr_bits-8{1'b0}}, next_instruction_value.opcode}) :
            next_instruction_address;
    else
        next_addr = current.next;
end

always @(posedge clk)
    addr <= next_addr;

always @(posedge clk)
    current <= mem[next_addr];

always_ff @(posedge clk)
    if (fifo_rd_en)
        cur_instruction <= next_instruction_value;

`ifdef verilator
export "DPI-C" function get_microcode_address;

function bit [addr_bits-1:0] get_microcode_address;
    get_microcode_address = addr;
endfunction

export "DPI-C" function get_ext_int_yield;

function bit get_ext_int_yield;
    get_ext_int_yield = current.ext_int_yield;
endfunction

int microcode_coverage[num_instructions];

always_ff @(posedge clk)
    microcode_coverage[addr] <= microcode_coverage[addr] + 1;

export "DPI-C" function get_microcode_num_instructions;

function int get_microcode_num_instructions;
    get_microcode_num_instructions = num_instructions;
endfunction

export "DPI-C" function get_microcode_coverage_bin;

function int get_microcode_coverage_bin;
    input int bin;
    get_microcode_coverage_bin = microcode_coverage[bin];
endfunction
`endif

endmodule